magic
tech sky130A
magscale 1 2
timestamp 1635531245
<< locali >>
rect 190377 57443 190411 57749
rect 190929 57103 190963 57477
rect 221841 57035 221875 57409
rect 248337 57035 248371 57409
rect 384405 57171 384439 57477
rect 394709 57171 394743 57409
rect 349905 5763 349939 5865
rect 350089 5627 350123 5797
rect 391949 5627 391983 6137
rect 398021 5559 398055 6137
rect 398113 5559 398147 6205
rect 164801 3587 164835 3893
rect 452485 3655 452519 3689
rect 452485 3621 452761 3655
rect 454417 3587 454451 4165
rect 452519 3553 452853 3587
rect 277225 3383 277259 3553
rect 461041 3383 461075 4029
rect 461225 3859 461259 3961
rect 515689 3791 515723 3893
rect 461501 3451 461535 3689
rect 487169 3519 487203 3689
rect 513791 3281 514033 3315
rect 514125 3179 514159 3689
rect 515781 3587 515815 3893
<< viali >>
rect 190377 57749 190411 57783
rect 190377 57409 190411 57443
rect 190929 57477 190963 57511
rect 384405 57477 384439 57511
rect 190929 57069 190963 57103
rect 221841 57409 221875 57443
rect 221841 57001 221875 57035
rect 248337 57409 248371 57443
rect 384405 57137 384439 57171
rect 394709 57409 394743 57443
rect 394709 57137 394743 57171
rect 248337 57001 248371 57035
rect 398113 6205 398147 6239
rect 391949 6137 391983 6171
rect 349905 5865 349939 5899
rect 349905 5729 349939 5763
rect 350089 5797 350123 5831
rect 350089 5593 350123 5627
rect 391949 5593 391983 5627
rect 398021 6137 398055 6171
rect 398021 5525 398055 5559
rect 398113 5525 398147 5559
rect 454417 4165 454451 4199
rect 164801 3893 164835 3927
rect 452485 3689 452519 3723
rect 452761 3621 452795 3655
rect 164801 3553 164835 3587
rect 277225 3553 277259 3587
rect 452485 3553 452519 3587
rect 452853 3553 452887 3587
rect 454417 3553 454451 3587
rect 461041 4029 461075 4063
rect 277225 3349 277259 3383
rect 461225 3961 461259 3995
rect 461225 3825 461259 3859
rect 515689 3893 515723 3927
rect 515689 3757 515723 3791
rect 515781 3893 515815 3927
rect 461501 3689 461535 3723
rect 487169 3689 487203 3723
rect 487169 3485 487203 3519
rect 514125 3689 514159 3723
rect 461501 3417 461535 3451
rect 461041 3349 461075 3383
rect 513757 3281 513791 3315
rect 514033 3281 514067 3315
rect 515781 3553 515815 3587
rect 514125 3145 514159 3179
<< metal1 >>
rect 430482 700408 430488 700460
rect 430540 700448 430546 700460
rect 462314 700448 462320 700460
rect 430540 700420 462320 700448
rect 430540 700408 430546 700420
rect 462314 700408 462320 700420
rect 462372 700408 462378 700460
rect 482922 700408 482928 700460
rect 482980 700448 482986 700460
rect 527174 700448 527180 700460
rect 482980 700420 527180 700448
rect 482980 700408 482986 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 393222 700340 393228 700392
rect 393280 700380 393286 700392
rect 413646 700380 413652 700392
rect 393280 700352 413652 700380
rect 393280 700340 393286 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 444282 700340 444288 700392
rect 444340 700380 444346 700392
rect 478506 700380 478512 700392
rect 444340 700352 478512 700380
rect 444340 700340 444346 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 495342 700340 495348 700392
rect 495400 700380 495406 700392
rect 543458 700380 543464 700392
rect 495400 700352 543464 700380
rect 495400 700340 495406 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 340782 700272 340788 700324
rect 340840 700312 340846 700324
rect 348786 700312 348792 700324
rect 340840 700284 348792 700312
rect 340840 700272 340846 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 354582 700272 354588 700324
rect 354640 700312 354646 700324
rect 364978 700312 364984 700324
rect 354640 700284 364984 700312
rect 354640 700272 354646 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 379422 700272 379428 700324
rect 379480 700312 379486 700324
rect 397454 700312 397460 700324
rect 379480 700284 397460 700312
rect 379480 700272 379486 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 405642 700272 405648 700324
rect 405700 700312 405706 700324
rect 429838 700312 429844 700324
rect 405700 700284 429844 700312
rect 405700 700272 405706 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 456702 700272 456708 700324
rect 456760 700312 456766 700324
rect 494790 700312 494796 700324
rect 456760 700284 494796 700312
rect 456760 700272 456766 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 507762 700272 507768 700324
rect 507820 700312 507826 700324
rect 559650 700312 559656 700324
rect 507820 700284 559656 700312
rect 507820 700272 507826 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 328362 699660 328368 699712
rect 328420 699700 328426 699712
rect 332502 699700 332508 699712
rect 328420 699672 332508 699700
rect 328420 699660 328426 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 522298 696940 522304 696992
rect 522356 696980 522362 696992
rect 580166 696980 580172 696992
rect 522356 696952 580172 696980
rect 522356 696940 522362 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 522390 683136 522396 683188
rect 522448 683176 522454 683188
rect 580166 683176 580172 683188
rect 522448 683148 580172 683176
rect 522448 683136 522454 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 522482 670692 522488 670744
rect 522540 670732 522546 670744
rect 580166 670732 580172 670744
rect 522540 670704 580172 670732
rect 522540 670692 522546 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 300762 655460 300768 655512
rect 300820 655500 300826 655512
rect 302326 655500 302332 655512
rect 300820 655472 302332 655500
rect 300820 655460 300826 655472
rect 302326 655460 302332 655472
rect 302384 655460 302390 655512
rect 353570 655460 353576 655512
rect 353628 655500 353634 655512
rect 354582 655500 354588 655512
rect 353628 655472 354588 655500
rect 353628 655460 353634 655472
rect 354582 655460 354588 655472
rect 354640 655460 354646 655512
rect 443178 655460 443184 655512
rect 443236 655500 443242 655512
rect 444282 655500 444288 655512
rect 443236 655472 444288 655500
rect 443236 655460 443242 655472
rect 444282 655460 444288 655472
rect 444340 655460 444346 655512
rect 455966 655460 455972 655512
rect 456024 655500 456030 655512
rect 456702 655500 456708 655512
rect 456024 655472 456708 655500
rect 456024 655460 456030 655472
rect 456702 655460 456708 655472
rect 456760 655460 456766 655512
rect 481634 655460 481640 655512
rect 481692 655500 481698 655512
rect 482922 655500 482928 655512
rect 481692 655472 482928 655500
rect 481692 655460 481698 655472
rect 482922 655460 482928 655472
rect 482980 655460 482986 655512
rect 494422 654984 494428 655036
rect 494480 655024 494486 655036
rect 495342 655024 495348 655036
rect 494480 654996 495348 655024
rect 494480 654984 494486 654996
rect 495342 654984 495348 654996
rect 495400 654984 495406 655036
rect 41322 654916 41328 654968
rect 41380 654956 41386 654968
rect 97534 654956 97540 654968
rect 41380 654928 97540 654956
rect 41380 654916 41386 654928
rect 97534 654916 97540 654928
rect 97592 654916 97598 654968
rect 106182 654916 106188 654968
rect 106240 654956 106246 654968
rect 148778 654956 148784 654968
rect 106240 654928 148784 654956
rect 106240 654916 106246 654928
rect 148778 654916 148784 654928
rect 148836 654916 148842 654968
rect 171042 654916 171048 654968
rect 171100 654956 171106 654968
rect 199930 654956 199936 654968
rect 171100 654928 199936 654956
rect 171100 654916 171106 654928
rect 199930 654916 199936 654928
rect 199988 654916 199994 654968
rect 24762 654848 24768 654900
rect 24820 654888 24826 654900
rect 84746 654888 84752 654900
rect 24820 654860 84752 654888
rect 24820 654848 24826 654860
rect 84746 654848 84752 654860
rect 84804 654848 84810 654900
rect 89622 654848 89628 654900
rect 89680 654888 89686 654900
rect 135990 654888 135996 654900
rect 89680 654860 135996 654888
rect 89680 654848 89686 654860
rect 135990 654848 135996 654860
rect 136048 654848 136054 654900
rect 154482 654848 154488 654900
rect 154540 654888 154546 654900
rect 187142 654888 187148 654900
rect 154540 654860 187148 654888
rect 154540 654848 154546 654860
rect 187142 654848 187148 654860
rect 187200 654848 187206 654900
rect 219342 654848 219348 654900
rect 219400 654888 219406 654900
rect 238294 654888 238300 654900
rect 219400 654860 238300 654888
rect 219400 654848 219406 654860
rect 238294 654848 238300 654860
rect 238352 654848 238358 654900
rect 8202 654780 8208 654832
rect 8260 654820 8266 654832
rect 72970 654820 72976 654832
rect 8260 654792 72976 654820
rect 8260 654780 8266 654792
rect 72970 654780 72976 654792
rect 73028 654780 73034 654832
rect 73062 654780 73068 654832
rect 73120 654820 73126 654832
rect 123110 654820 123116 654832
rect 73120 654792 123116 654820
rect 73120 654780 73126 654792
rect 123110 654780 123116 654792
rect 123168 654780 123174 654832
rect 137922 654780 137928 654832
rect 137980 654820 137986 654832
rect 174354 654820 174360 654832
rect 137980 654792 174360 654820
rect 137980 654780 137986 654792
rect 174354 654780 174360 654792
rect 174412 654780 174418 654832
rect 202782 654780 202788 654832
rect 202840 654820 202846 654832
rect 225506 654820 225512 654832
rect 202840 654792 225512 654820
rect 202840 654780 202846 654792
rect 225506 654780 225512 654792
rect 225564 654780 225570 654832
rect 235902 654780 235908 654832
rect 235960 654820 235966 654832
rect 251174 654820 251180 654832
rect 235960 654792 251180 654820
rect 235960 654780 235966 654792
rect 251174 654780 251180 654792
rect 251232 654780 251238 654832
rect 267642 654780 267648 654832
rect 267700 654820 267706 654832
rect 276750 654820 276756 654832
rect 267700 654792 276756 654820
rect 267700 654780 267706 654792
rect 276750 654780 276756 654792
rect 276808 654780 276814 654832
rect 404814 654780 404820 654832
rect 404872 654820 404878 654832
rect 405642 654820 405648 654832
rect 404872 654792 405648 654820
rect 404872 654780 404878 654792
rect 405642 654780 405648 654792
rect 405700 654780 405706 654832
rect 392026 654576 392032 654628
rect 392084 654616 392090 654628
rect 393222 654616 393228 654628
rect 392084 654588 393228 654616
rect 392084 654576 392090 654588
rect 393222 654576 393228 654588
rect 393280 654576 393286 654628
rect 284202 654372 284208 654424
rect 284260 654412 284266 654424
rect 289538 654412 289544 654424
rect 284260 654384 289544 654412
rect 284260 654372 284266 654384
rect 289538 654372 289544 654384
rect 289596 654372 289602 654424
rect 507210 654372 507216 654424
rect 507268 654412 507274 654424
rect 507762 654412 507768 654424
rect 507268 654384 507768 654412
rect 507268 654372 507274 654384
rect 507762 654372 507768 654384
rect 507820 654372 507826 654424
rect 522298 643084 522304 643136
rect 522356 643124 522362 643136
rect 580166 643124 580172 643136
rect 522356 643096 580172 643124
rect 522356 643084 522362 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 641656 3424 641708
rect 3476 641696 3482 641708
rect 69014 641696 69020 641708
rect 3476 641668 69020 641696
rect 3476 641656 3482 641668
rect 69014 641656 69020 641668
rect 69072 641656 69078 641708
rect 522390 630640 522396 630692
rect 522448 630680 522454 630692
rect 580166 630680 580172 630692
rect 522448 630652 580172 630680
rect 522448 630640 522454 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 630572 3516 630624
rect 3568 630612 3574 630624
rect 69014 630612 69020 630624
rect 3568 630584 69020 630612
rect 3568 630572 3574 630584
rect 69014 630572 69020 630584
rect 69072 630572 69078 630624
rect 3602 619556 3608 619608
rect 3660 619596 3666 619608
rect 69014 619596 69020 619608
rect 3660 619568 69020 619596
rect 3660 619556 3666 619568
rect 69014 619556 69020 619568
rect 69072 619556 69078 619608
rect 522482 616836 522488 616888
rect 522540 616876 522546 616888
rect 580166 616876 580172 616888
rect 522540 616848 580172 616876
rect 522540 616836 522546 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 597456 3424 597508
rect 3476 597496 3482 597508
rect 69014 597496 69020 597508
rect 3476 597468 69020 597496
rect 3476 597456 3482 597468
rect 69014 597456 69020 597468
rect 69072 597456 69078 597508
rect 522298 590656 522304 590708
rect 522356 590696 522362 590708
rect 579798 590696 579804 590708
rect 522356 590668 579804 590696
rect 522356 590656 522362 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3510 585080 3516 585132
rect 3568 585120 3574 585132
rect 69014 585120 69020 585132
rect 3568 585092 69020 585120
rect 3568 585080 3574 585092
rect 69014 585080 69020 585092
rect 69072 585080 69078 585132
rect 522390 576852 522396 576904
rect 522448 576892 522454 576904
rect 580166 576892 580172 576904
rect 522448 576864 580172 576892
rect 522448 576852 522454 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3602 573996 3608 574048
rect 3660 574036 3666 574048
rect 69014 574036 69020 574048
rect 3660 574008 69020 574036
rect 3660 573996 3666 574008
rect 69014 573996 69020 574008
rect 69072 573996 69078 574048
rect 522482 563048 522488 563100
rect 522540 563088 522546 563100
rect 579798 563088 579804 563100
rect 522540 563060 579804 563088
rect 522540 563048 522546 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 551964 3424 552016
rect 3476 552004 3482 552016
rect 69014 552004 69020 552016
rect 3476 551976 69020 552004
rect 3476 551964 3482 551976
rect 69014 551964 69020 551976
rect 69072 551964 69078 552016
rect 3510 540880 3516 540932
rect 3568 540920 3574 540932
rect 69014 540920 69020 540932
rect 3568 540892 69020 540920
rect 3568 540880 3574 540892
rect 69014 540880 69020 540892
rect 69072 540880 69078 540932
rect 522298 536800 522304 536852
rect 522356 536840 522362 536852
rect 580166 536840 580172 536852
rect 522356 536812 580172 536840
rect 522356 536800 522362 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3602 529864 3608 529916
rect 3660 529904 3666 529916
rect 69014 529904 69020 529916
rect 3660 529876 69020 529904
rect 3660 529864 3666 529876
rect 69014 529864 69020 529876
rect 69072 529864 69078 529916
rect 522390 524424 522396 524476
rect 522448 524464 522454 524476
rect 580166 524464 580172 524476
rect 522448 524436 580172 524464
rect 522448 524424 522454 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 522298 510620 522304 510672
rect 522356 510660 522362 510672
rect 580166 510660 580172 510672
rect 522356 510632 580172 510660
rect 522356 510620 522362 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3418 507764 3424 507816
rect 3476 507804 3482 507816
rect 69014 507804 69020 507816
rect 3476 507776 69020 507804
rect 3476 507764 3482 507776
rect 69014 507764 69020 507776
rect 69072 507764 69078 507816
rect 3510 496748 3516 496800
rect 3568 496788 3574 496800
rect 69014 496788 69020 496800
rect 3568 496760 69020 496788
rect 3568 496748 3574 496760
rect 69014 496748 69020 496760
rect 69072 496748 69078 496800
rect 3418 485732 3424 485784
rect 3476 485772 3482 485784
rect 69014 485772 69020 485784
rect 3476 485744 69020 485772
rect 3476 485732 3482 485744
rect 69014 485732 69020 485744
rect 69072 485732 69078 485784
rect 522298 484372 522304 484424
rect 522356 484412 522362 484424
rect 580166 484412 580172 484424
rect 522356 484384 580172 484412
rect 522356 484372 522362 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 522390 470568 522396 470620
rect 522448 470608 522454 470620
rect 579982 470608 579988 470620
rect 522448 470580 579988 470608
rect 522448 470568 522454 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3418 462272 3424 462324
rect 3476 462312 3482 462324
rect 69014 462312 69020 462324
rect 3476 462284 69020 462312
rect 3476 462272 3482 462284
rect 69014 462272 69020 462284
rect 69072 462272 69078 462324
rect 522298 456764 522304 456816
rect 522356 456804 522362 456816
rect 580166 456804 580172 456816
rect 522356 456776 580172 456804
rect 522356 456764 522362 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3510 451188 3516 451240
rect 3568 451228 3574 451240
rect 69014 451228 69020 451240
rect 3568 451200 69020 451228
rect 3568 451188 3574 451200
rect 69014 451188 69020 451200
rect 69072 451188 69078 451240
rect 3418 440172 3424 440224
rect 3476 440212 3482 440224
rect 69014 440212 69020 440224
rect 3476 440184 69020 440212
rect 3476 440172 3482 440184
rect 69014 440172 69020 440184
rect 69072 440172 69078 440224
rect 522942 430584 522948 430636
rect 523000 430624 523006 430636
rect 580166 430624 580172 430636
rect 523000 430596 580172 430624
rect 523000 430584 523006 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 522942 418140 522948 418192
rect 523000 418180 523006 418192
rect 580166 418180 580172 418192
rect 523000 418152 580172 418180
rect 523000 418140 523006 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 418072 3332 418124
rect 3384 418112 3390 418124
rect 69014 418112 69020 418124
rect 3384 418084 69020 418112
rect 3384 418072 3390 418084
rect 69014 418072 69020 418084
rect 69072 418072 69078 418124
rect 3418 407056 3424 407108
rect 3476 407096 3482 407108
rect 69014 407096 69020 407108
rect 3476 407068 69020 407096
rect 3476 407056 3482 407068
rect 69014 407056 69020 407068
rect 69072 407056 69078 407108
rect 522022 404336 522028 404388
rect 522080 404376 522086 404388
rect 580166 404376 580172 404388
rect 522080 404348 580172 404376
rect 522080 404336 522086 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 2866 395972 2872 396024
rect 2924 396012 2930 396024
rect 69014 396012 69020 396024
rect 2924 395984 69020 396012
rect 2924 395972 2930 395984
rect 69014 395972 69020 395984
rect 69072 395972 69078 396024
rect 522942 378768 522948 378820
rect 523000 378808 523006 378820
rect 580166 378808 580172 378820
rect 523000 378780 580172 378808
rect 523000 378768 523006 378780
rect 580166 378768 580172 378780
rect 580224 378768 580230 378820
rect 3418 372580 3424 372632
rect 3476 372620 3482 372632
rect 69014 372620 69020 372632
rect 3476 372592 69020 372620
rect 3476 372580 3482 372592
rect 69014 372580 69020 372592
rect 69072 372580 69078 372632
rect 522942 365644 522948 365696
rect 523000 365684 523006 365696
rect 580166 365684 580172 365696
rect 523000 365656 580172 365684
rect 523000 365644 523006 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3418 361564 3424 361616
rect 3476 361604 3482 361616
rect 69014 361604 69020 361616
rect 3476 361576 69020 361604
rect 3476 361564 3482 361576
rect 69014 361564 69020 361576
rect 69072 361564 69078 361616
rect 522942 353200 522948 353252
rect 523000 353240 523006 353252
rect 580166 353240 580172 353252
rect 523000 353212 580172 353240
rect 523000 353200 523006 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 2866 349120 2872 349172
rect 2924 349160 2930 349172
rect 69014 349160 69020 349172
rect 2924 349132 69020 349160
rect 2924 349120 2930 349132
rect 69014 349120 69020 349132
rect 69072 349120 69078 349172
rect 2866 327088 2872 327140
rect 2924 327128 2930 327140
rect 69014 327128 69020 327140
rect 2924 327100 69020 327128
rect 2924 327088 2930 327100
rect 69014 327088 69020 327100
rect 69072 327088 69078 327140
rect 522298 325592 522304 325644
rect 522356 325632 522362 325644
rect 580166 325632 580172 325644
rect 522356 325604 580172 325632
rect 522356 325592 522362 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3510 316004 3516 316056
rect 3568 316044 3574 316056
rect 69014 316044 69020 316056
rect 3568 316016 69020 316044
rect 3568 316004 3574 316016
rect 69014 316004 69020 316016
rect 69072 316004 69078 316056
rect 522298 313216 522304 313268
rect 522356 313256 522362 313268
rect 580166 313256 580172 313268
rect 522356 313228 580172 313256
rect 522356 313216 522362 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 69014 305028 69020 305040
rect 3476 305000 69020 305028
rect 3476 304988 3482 305000
rect 69014 304988 69020 305000
rect 69072 304988 69078 305040
rect 522298 299412 522304 299464
rect 522356 299452 522362 299464
rect 580166 299452 580172 299464
rect 522356 299424 580172 299452
rect 522356 299412 522362 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3418 282888 3424 282940
rect 3476 282928 3482 282940
rect 69014 282928 69020 282940
rect 3476 282900 69020 282928
rect 3476 282888 3482 282900
rect 69014 282888 69020 282900
rect 69072 282888 69078 282940
rect 522390 273164 522396 273216
rect 522448 273204 522454 273216
rect 580166 273204 580172 273216
rect 522448 273176 580172 273204
rect 522448 273164 522454 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3510 271872 3516 271924
rect 3568 271912 3574 271924
rect 69014 271912 69020 271924
rect 3568 271884 69020 271912
rect 3568 271872 3574 271884
rect 69014 271872 69020 271884
rect 69072 271872 69078 271924
rect 3418 260856 3424 260908
rect 3476 260896 3482 260908
rect 69014 260896 69020 260908
rect 3476 260868 69020 260896
rect 3476 260856 3482 260868
rect 69014 260856 69020 260868
rect 69072 260856 69078 260908
rect 522298 259360 522304 259412
rect 522356 259400 522362 259412
rect 580166 259400 580172 259412
rect 522356 259372 580172 259400
rect 522356 259360 522362 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 522390 245556 522396 245608
rect 522448 245596 522454 245608
rect 580166 245596 580172 245608
rect 522448 245568 580172 245596
rect 522448 245556 522454 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 238756 3516 238808
rect 3568 238796 3574 238808
rect 69014 238796 69020 238808
rect 3568 238768 69020 238796
rect 3568 238756 3574 238768
rect 69014 238756 69020 238768
rect 69072 238756 69078 238808
rect 522298 233180 522304 233232
rect 522356 233220 522362 233232
rect 579982 233220 579988 233232
rect 522356 233192 579988 233220
rect 522356 233180 522362 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3602 226312 3608 226364
rect 3660 226352 3666 226364
rect 69014 226352 69020 226364
rect 3660 226324 69020 226352
rect 3660 226312 3666 226324
rect 69014 226312 69020 226324
rect 69072 226312 69078 226364
rect 522390 219376 522396 219428
rect 522448 219416 522454 219428
rect 580166 219416 580172 219428
rect 522448 219388 580172 219416
rect 522448 219376 522454 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3418 215296 3424 215348
rect 3476 215336 3482 215348
rect 69014 215336 69020 215348
rect 3476 215308 69020 215336
rect 3476 215296 3482 215308
rect 69014 215296 69020 215308
rect 69072 215296 69078 215348
rect 522298 206932 522304 206984
rect 522356 206972 522362 206984
rect 579798 206972 579804 206984
rect 522356 206944 579804 206972
rect 522356 206932 522362 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3602 193196 3608 193248
rect 3660 193236 3666 193248
rect 69014 193236 69020 193248
rect 3660 193208 69020 193236
rect 3660 193196 3666 193208
rect 69014 193196 69020 193208
rect 69072 193196 69078 193248
rect 522482 193128 522488 193180
rect 522540 193168 522546 193180
rect 580166 193168 580172 193180
rect 522540 193140 580172 193168
rect 522540 193128 522546 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 182180 3516 182232
rect 3568 182220 3574 182232
rect 69014 182220 69020 182232
rect 3568 182192 69020 182220
rect 3568 182180 3574 182192
rect 69014 182180 69020 182192
rect 69072 182180 69078 182232
rect 522390 179324 522396 179376
rect 522448 179364 522454 179376
rect 580166 179364 580172 179376
rect 522448 179336 580172 179364
rect 522448 179324 522454 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 3418 171096 3424 171148
rect 3476 171136 3482 171148
rect 69014 171136 69020 171148
rect 3476 171108 69020 171136
rect 3476 171096 3482 171108
rect 69014 171096 69020 171108
rect 69072 171096 69078 171148
rect 522298 166948 522304 167000
rect 522356 166988 522362 167000
rect 580166 166988 580172 167000
rect 522356 166960 580172 166988
rect 522356 166948 522362 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 522482 153144 522488 153196
rect 522540 153184 522546 153196
rect 580166 153184 580172 153196
rect 522540 153156 580172 153184
rect 522540 153144 522546 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3694 149064 3700 149116
rect 3752 149104 3758 149116
rect 69014 149104 69020 149116
rect 3752 149076 69020 149104
rect 3752 149064 3758 149076
rect 69014 149064 69020 149076
rect 69072 149064 69078 149116
rect 522390 139340 522396 139392
rect 522448 139380 522454 139392
rect 580166 139380 580172 139392
rect 522448 139352 580172 139380
rect 522448 139340 522454 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3602 137980 3608 138032
rect 3660 138020 3666 138032
rect 69014 138020 69020 138032
rect 3660 137992 69020 138020
rect 3660 137980 3666 137992
rect 69014 137980 69020 137992
rect 69072 137980 69078 138032
rect 3510 126964 3516 127016
rect 3568 127004 3574 127016
rect 69014 127004 69020 127016
rect 3568 126976 69020 127004
rect 3568 126964 3574 126976
rect 69014 126964 69020 126976
rect 69072 126964 69078 127016
rect 522298 126896 522304 126948
rect 522356 126936 522362 126948
rect 580166 126936 580172 126948
rect 522356 126908 580172 126936
rect 522356 126896 522362 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3418 114520 3424 114572
rect 3476 114560 3482 114572
rect 69014 114560 69020 114572
rect 3476 114532 69020 114560
rect 3476 114520 3482 114532
rect 69014 114520 69020 114532
rect 69072 114520 69078 114572
rect 522574 113092 522580 113144
rect 522632 113132 522638 113144
rect 579798 113132 579804 113144
rect 522632 113104 579804 113132
rect 522632 113092 522638 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3786 103504 3792 103556
rect 3844 103544 3850 103556
rect 69014 103544 69020 103556
rect 3844 103516 69020 103544
rect 3844 103504 3850 103516
rect 69014 103504 69020 103516
rect 69072 103504 69078 103556
rect 522482 100648 522488 100700
rect 522540 100688 522546 100700
rect 580166 100688 580172 100700
rect 522540 100660 580172 100688
rect 522540 100648 522546 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3694 92488 3700 92540
rect 3752 92528 3758 92540
rect 69014 92528 69020 92540
rect 3752 92500 69020 92528
rect 3752 92488 3758 92500
rect 69014 92488 69020 92500
rect 69072 92488 69078 92540
rect 522390 86912 522396 86964
rect 522448 86952 522454 86964
rect 580166 86952 580172 86964
rect 522448 86924 580172 86952
rect 522448 86912 522454 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3602 81404 3608 81456
rect 3660 81444 3666 81456
rect 69014 81444 69020 81456
rect 3660 81416 69020 81444
rect 3660 81404 3666 81416
rect 69014 81404 69020 81416
rect 69072 81404 69078 81456
rect 522298 73108 522304 73160
rect 522356 73148 522362 73160
rect 580166 73148 580172 73160
rect 522356 73120 580172 73148
rect 522356 73108 522362 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 70388 3516 70440
rect 3568 70428 3574 70440
rect 69014 70428 69020 70440
rect 3568 70400 69020 70428
rect 3568 70388 3574 70400
rect 69014 70388 69020 70400
rect 69072 70388 69078 70440
rect 3418 60732 3424 60784
rect 3476 60772 3482 60784
rect 69014 60772 69020 60784
rect 3476 60744 69020 60772
rect 3476 60732 3482 60744
rect 69014 60732 69020 60744
rect 69072 60732 69078 60784
rect 522666 60664 522672 60716
rect 522724 60704 522730 60716
rect 580166 60704 580172 60716
rect 522724 60676 580172 60704
rect 522724 60664 522730 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 295334 59780 295340 59832
rect 295392 59820 295398 59832
rect 296310 59820 296316 59832
rect 295392 59792 296316 59820
rect 295392 59780 295398 59792
rect 296310 59780 296316 59792
rect 296368 59780 296374 59832
rect 313366 59780 313372 59832
rect 313424 59820 313430 59832
rect 314526 59820 314532 59832
rect 313424 59792 314532 59820
rect 313424 59780 313430 59792
rect 314526 59780 314532 59792
rect 314584 59780 314590 59832
rect 324314 59780 324320 59832
rect 324372 59820 324378 59832
rect 325382 59820 325388 59832
rect 324372 59792 325388 59820
rect 324372 59780 324378 59792
rect 325382 59780 325388 59792
rect 325440 59780 325446 59832
rect 427814 59780 427820 59832
rect 427872 59820 427878 59832
rect 428974 59820 428980 59832
rect 427872 59792 428980 59820
rect 427872 59780 427878 59792
rect 428974 59780 428980 59792
rect 429032 59780 429038 59832
rect 430574 59780 430580 59832
rect 430632 59820 430638 59832
rect 431734 59820 431740 59832
rect 430632 59792 431740 59820
rect 430632 59780 430638 59792
rect 431734 59780 431740 59792
rect 431792 59780 431798 59832
rect 436094 59780 436100 59832
rect 436152 59820 436158 59832
rect 437162 59820 437168 59832
rect 436152 59792 437168 59820
rect 436152 59780 436158 59792
rect 437162 59780 437168 59792
rect 437220 59780 437226 59832
rect 438854 59780 438860 59832
rect 438912 59820 438918 59832
rect 439922 59820 439928 59832
rect 438912 59792 439928 59820
rect 438912 59780 438918 59792
rect 439922 59780 439928 59792
rect 439980 59780 439986 59832
rect 456794 59780 456800 59832
rect 456852 59820 456858 59832
rect 458046 59820 458052 59832
rect 456852 59792 458052 59820
rect 456852 59780 456858 59792
rect 458046 59780 458052 59792
rect 458104 59780 458110 59832
rect 467834 59780 467840 59832
rect 467892 59820 467898 59832
rect 468994 59820 469000 59832
rect 467892 59792 469000 59820
rect 467892 59780 467898 59792
rect 468994 59780 469000 59792
rect 469052 59780 469058 59832
rect 155862 57876 155868 57928
rect 155920 57916 155926 57928
rect 291746 57916 291752 57928
rect 155920 57888 291752 57916
rect 155920 57876 155926 57888
rect 291746 57876 291752 57888
rect 291804 57876 291810 57928
rect 383654 57876 383660 57928
rect 383712 57916 383718 57928
rect 384850 57916 384856 57928
rect 383712 57888 384856 57916
rect 383712 57876 383718 57888
rect 384850 57876 384856 57888
rect 384908 57876 384914 57928
rect 469122 57876 469128 57928
rect 469180 57916 469186 57928
rect 487982 57916 487988 57928
rect 469180 57888 487988 57916
rect 469180 57876 469186 57888
rect 487982 57876 487988 57888
rect 488040 57876 488046 57928
rect 153102 57808 153108 57860
rect 153160 57848 153166 57860
rect 290826 57848 290832 57860
rect 153160 57820 290832 57848
rect 153160 57808 153166 57820
rect 290826 57808 290832 57820
rect 290884 57808 290890 57860
rect 375466 57808 375472 57860
rect 375524 57848 375530 57860
rect 443638 57848 443644 57860
rect 375524 57820 443644 57848
rect 375524 57808 375530 57820
rect 443638 57808 443644 57820
rect 443696 57808 443702 57860
rect 473262 57808 473268 57860
rect 473320 57848 473326 57860
rect 488902 57848 488908 57860
rect 473320 57820 488908 57848
rect 473320 57808 473326 57820
rect 488902 57808 488908 57820
rect 488960 57808 488966 57860
rect 136542 57740 136548 57792
rect 136600 57780 136606 57792
rect 170858 57780 170864 57792
rect 136600 57752 170864 57780
rect 136600 57740 136606 57752
rect 170858 57740 170864 57752
rect 170916 57740 170922 57792
rect 184658 57740 184664 57792
rect 184716 57780 184722 57792
rect 186958 57780 186964 57792
rect 184716 57752 186964 57780
rect 184716 57740 184722 57752
rect 186958 57740 186964 57752
rect 187016 57740 187022 57792
rect 187326 57740 187332 57792
rect 187384 57780 187390 57792
rect 190365 57783 190423 57789
rect 190365 57780 190377 57783
rect 187384 57752 190377 57780
rect 187384 57740 187390 57752
rect 190365 57749 190377 57752
rect 190411 57749 190423 57783
rect 190365 57743 190423 57749
rect 200114 57740 200120 57792
rect 200172 57780 200178 57792
rect 201310 57780 201316 57792
rect 200172 57752 201316 57780
rect 200172 57740 200178 57752
rect 201310 57740 201316 57752
rect 201368 57740 201374 57792
rect 218238 57740 218244 57792
rect 218296 57780 218302 57792
rect 222838 57780 222844 57792
rect 218296 57752 222844 57780
rect 218296 57740 218302 57752
rect 222838 57740 222844 57752
rect 222896 57740 222902 57792
rect 225506 57740 225512 57792
rect 225564 57780 225570 57792
rect 233878 57780 233884 57792
rect 225564 57752 233884 57780
rect 225564 57740 225570 57752
rect 233878 57740 233884 57752
rect 233936 57740 233942 57792
rect 234614 57740 234620 57792
rect 234672 57780 234678 57792
rect 374638 57780 374644 57792
rect 234672 57752 374644 57780
rect 234672 57740 234678 57752
rect 374638 57740 374644 57752
rect 374696 57740 374702 57792
rect 380894 57740 380900 57792
rect 380952 57780 380958 57792
rect 449158 57780 449164 57792
rect 380952 57752 449164 57780
rect 380952 57740 380958 57752
rect 449158 57740 449164 57752
rect 449216 57740 449222 57792
rect 466362 57740 466368 57792
rect 466420 57780 466426 57792
rect 487154 57780 487160 57792
rect 466420 57752 487160 57780
rect 466420 57740 466426 57752
rect 487154 57740 487160 57752
rect 487212 57740 487218 57792
rect 148962 57672 148968 57724
rect 149020 57712 149026 57724
rect 289906 57712 289912 57724
rect 149020 57684 289912 57712
rect 149020 57672 149026 57684
rect 289906 57672 289912 57684
rect 289964 57672 289970 57724
rect 377398 57672 377404 57724
rect 377456 57712 377462 57724
rect 455414 57712 455420 57724
rect 377456 57684 455420 57712
rect 377456 57672 377462 57684
rect 455414 57672 455420 57684
rect 455472 57672 455478 57724
rect 462222 57672 462228 57724
rect 462280 57712 462286 57724
rect 486234 57712 486240 57724
rect 462280 57684 486240 57712
rect 462280 57672 462286 57684
rect 486234 57672 486240 57684
rect 486292 57672 486298 57724
rect 144822 57604 144828 57656
rect 144880 57644 144886 57656
rect 288986 57644 288992 57656
rect 144880 57616 288992 57644
rect 144880 57604 144886 57616
rect 288986 57604 288992 57616
rect 289044 57604 289050 57656
rect 305638 57604 305644 57656
rect 305696 57644 305702 57656
rect 321554 57644 321560 57656
rect 305696 57616 321560 57644
rect 305696 57604 305702 57616
rect 321554 57604 321560 57616
rect 321612 57604 321618 57656
rect 332594 57604 332600 57656
rect 332652 57644 332658 57656
rect 333514 57644 333520 57656
rect 332652 57616 333520 57644
rect 332652 57604 332658 57616
rect 333514 57604 333520 57616
rect 333572 57604 333578 57656
rect 335354 57604 335360 57656
rect 335412 57644 335418 57656
rect 336274 57644 336280 57656
rect 335412 57616 336280 57644
rect 335412 57604 335418 57616
rect 336274 57604 336280 57616
rect 336332 57604 336338 57656
rect 339954 57604 339960 57656
rect 340012 57644 340018 57656
rect 340782 57644 340788 57656
rect 340012 57616 340788 57644
rect 340012 57604 340018 57616
rect 340782 57604 340788 57616
rect 340840 57604 340846 57656
rect 340874 57604 340880 57656
rect 340932 57644 340938 57656
rect 342070 57644 342076 57656
rect 340932 57616 342076 57644
rect 340932 57604 340938 57616
rect 342070 57604 342076 57616
rect 342128 57604 342134 57656
rect 342714 57604 342720 57656
rect 342772 57644 342778 57656
rect 343542 57644 343548 57656
rect 342772 57616 343548 57644
rect 342772 57604 342778 57616
rect 343542 57604 343548 57616
rect 343600 57604 343606 57656
rect 343634 57604 343640 57656
rect 343692 57644 343698 57656
rect 344922 57644 344928 57656
rect 343692 57616 344928 57644
rect 343692 57604 343698 57616
rect 344922 57604 344928 57616
rect 344980 57604 344986 57656
rect 345474 57604 345480 57656
rect 345532 57644 345538 57656
rect 346302 57644 346308 57656
rect 345532 57616 346308 57644
rect 345532 57604 345538 57616
rect 346302 57604 346308 57616
rect 346360 57604 346366 57656
rect 346394 57604 346400 57656
rect 346452 57644 346458 57656
rect 347590 57644 347596 57656
rect 346452 57616 347596 57644
rect 346452 57604 346458 57616
rect 347590 57604 347596 57616
rect 347648 57604 347654 57656
rect 348142 57604 348148 57656
rect 348200 57644 348206 57656
rect 348970 57644 348976 57656
rect 348200 57616 348976 57644
rect 348200 57604 348206 57616
rect 348970 57604 348976 57616
rect 349028 57604 349034 57656
rect 350902 57604 350908 57656
rect 350960 57644 350966 57656
rect 351730 57644 351736 57656
rect 350960 57616 351736 57644
rect 350960 57604 350966 57616
rect 351730 57604 351736 57616
rect 351788 57604 351794 57656
rect 353662 57604 353668 57656
rect 353720 57644 353726 57656
rect 354582 57644 354588 57656
rect 353720 57616 354588 57644
rect 353720 57604 353726 57616
rect 354582 57604 354588 57616
rect 354640 57604 354646 57656
rect 355410 57604 355416 57656
rect 355468 57644 355474 57656
rect 355962 57644 355968 57656
rect 355468 57616 355968 57644
rect 355468 57604 355474 57616
rect 355962 57604 355968 57616
rect 356020 57604 356026 57656
rect 356330 57604 356336 57656
rect 356388 57644 356394 57656
rect 357250 57644 357256 57656
rect 356388 57616 357256 57644
rect 356388 57604 356394 57616
rect 357250 57604 357256 57616
rect 357308 57604 357314 57656
rect 358170 57604 358176 57656
rect 358228 57644 358234 57656
rect 358722 57644 358728 57656
rect 358228 57616 358728 57644
rect 358228 57604 358234 57616
rect 358722 57604 358728 57616
rect 358780 57604 358786 57656
rect 359090 57604 359096 57656
rect 359148 57644 359154 57656
rect 360010 57644 360016 57656
rect 359148 57616 360016 57644
rect 359148 57604 359154 57616
rect 360010 57604 360016 57616
rect 360068 57604 360074 57656
rect 360930 57604 360936 57656
rect 360988 57644 360994 57656
rect 361482 57644 361488 57656
rect 360988 57616 361488 57644
rect 360988 57604 360994 57616
rect 361482 57604 361488 57616
rect 361540 57604 361546 57656
rect 363598 57604 363604 57656
rect 363656 57644 363662 57656
rect 364242 57644 364248 57656
rect 363656 57616 364248 57644
rect 363656 57604 363662 57616
rect 364242 57604 364248 57616
rect 364300 57604 364306 57656
rect 364518 57604 364524 57656
rect 364576 57644 364582 57656
rect 365530 57644 365536 57656
rect 364576 57616 365536 57644
rect 364576 57604 364582 57616
rect 365530 57604 365536 57616
rect 365588 57604 365594 57656
rect 366358 57604 366364 57656
rect 366416 57644 366422 57656
rect 367002 57644 367008 57656
rect 366416 57616 367008 57644
rect 366416 57604 366422 57616
rect 367002 57604 367008 57616
rect 367060 57604 367066 57656
rect 367278 57604 367284 57656
rect 367336 57644 367342 57656
rect 368382 57644 368388 57656
rect 367336 57616 368388 57644
rect 367336 57604 367342 57616
rect 368382 57604 368388 57616
rect 368440 57604 368446 57656
rect 369026 57604 369032 57656
rect 369084 57644 369090 57656
rect 369762 57644 369768 57656
rect 369084 57616 369768 57644
rect 369084 57604 369090 57616
rect 369762 57604 369768 57616
rect 369820 57604 369826 57656
rect 369946 57604 369952 57656
rect 370004 57644 370010 57656
rect 371050 57644 371056 57656
rect 370004 57616 371056 57644
rect 370004 57604 370010 57616
rect 371050 57604 371056 57616
rect 371108 57604 371114 57656
rect 371786 57604 371792 57656
rect 371844 57644 371850 57656
rect 372522 57644 372528 57656
rect 371844 57616 372528 57644
rect 371844 57604 371850 57616
rect 372522 57604 372528 57616
rect 372580 57604 372586 57656
rect 372706 57604 372712 57656
rect 372764 57644 372770 57656
rect 373810 57644 373816 57656
rect 372764 57616 373816 57644
rect 372764 57604 372770 57616
rect 373810 57604 373816 57616
rect 373868 57604 373874 57656
rect 374546 57604 374552 57656
rect 374604 57644 374610 57656
rect 375282 57644 375288 57656
rect 374604 57616 375288 57644
rect 374604 57604 374610 57616
rect 375282 57604 375288 57616
rect 375340 57604 375346 57656
rect 377214 57604 377220 57656
rect 377272 57644 377278 57656
rect 378042 57644 378048 57656
rect 377272 57616 378048 57644
rect 377272 57604 377278 57616
rect 378042 57604 378048 57616
rect 378100 57604 378106 57656
rect 378134 57604 378140 57656
rect 378192 57644 378198 57656
rect 379330 57644 379336 57656
rect 378192 57616 379336 57644
rect 378192 57604 378198 57616
rect 379330 57604 379336 57616
rect 379388 57604 379394 57656
rect 379974 57604 379980 57656
rect 380032 57644 380038 57656
rect 483658 57644 483664 57656
rect 380032 57616 483664 57644
rect 380032 57604 380038 57616
rect 483658 57604 483664 57616
rect 483716 57604 483722 57656
rect 496262 57604 496268 57656
rect 496320 57644 496326 57656
rect 497458 57644 497464 57656
rect 496320 57616 497464 57644
rect 496320 57604 496326 57616
rect 497458 57604 497464 57616
rect 497516 57604 497522 57656
rect 499022 57604 499028 57656
rect 499080 57644 499086 57656
rect 499482 57644 499488 57656
rect 499080 57616 499488 57644
rect 499080 57604 499086 57616
rect 499482 57604 499488 57616
rect 499540 57604 499546 57656
rect 499942 57604 499948 57656
rect 500000 57644 500006 57656
rect 500770 57644 500776 57656
rect 500000 57616 500776 57644
rect 500000 57604 500006 57616
rect 500770 57604 500776 57616
rect 500828 57604 500834 57656
rect 502610 57604 502616 57656
rect 502668 57644 502674 57656
rect 503622 57644 503628 57656
rect 502668 57616 503628 57644
rect 502668 57604 502674 57616
rect 503622 57604 503628 57616
rect 503680 57604 503686 57656
rect 505370 57604 505376 57656
rect 505428 57644 505434 57656
rect 506382 57644 506388 57656
rect 505428 57616 506388 57644
rect 505428 57604 505434 57616
rect 506382 57604 506388 57616
rect 506440 57604 506446 57656
rect 508130 57604 508136 57656
rect 508188 57644 508194 57656
rect 509050 57644 509056 57656
rect 508188 57616 509056 57644
rect 508188 57604 508194 57616
rect 509050 57604 509056 57616
rect 509108 57604 509114 57656
rect 509878 57604 509884 57656
rect 509936 57644 509942 57656
rect 510522 57644 510528 57656
rect 509936 57616 510528 57644
rect 509936 57604 509942 57616
rect 510522 57604 510528 57616
rect 510580 57604 510586 57656
rect 510798 57604 510804 57656
rect 510856 57644 510862 57656
rect 511810 57644 511816 57656
rect 510856 57616 511816 57644
rect 510856 57604 510862 57616
rect 511810 57604 511816 57616
rect 511868 57604 511874 57656
rect 512638 57604 512644 57656
rect 512696 57644 512702 57656
rect 513282 57644 513288 57656
rect 512696 57616 513288 57644
rect 512696 57604 512702 57616
rect 513282 57604 513288 57616
rect 513340 57604 513346 57656
rect 513558 57604 513564 57656
rect 513616 57644 513622 57656
rect 514662 57644 514668 57656
rect 513616 57616 514668 57644
rect 513616 57604 513622 57616
rect 514662 57604 514668 57616
rect 514720 57604 514726 57656
rect 515398 57604 515404 57656
rect 515456 57644 515462 57656
rect 516042 57644 516048 57656
rect 515456 57616 516048 57644
rect 515456 57604 515462 57616
rect 516042 57604 516048 57616
rect 516100 57604 516106 57656
rect 142062 57536 142068 57588
rect 142120 57576 142126 57588
rect 288158 57576 288164 57588
rect 142120 57548 288164 57576
rect 142120 57536 142126 57548
rect 288158 57536 288164 57548
rect 288216 57536 288222 57588
rect 288250 57536 288256 57588
rect 288308 57576 288314 57588
rect 300854 57576 300860 57588
rect 288308 57548 300860 57576
rect 288308 57536 288314 57548
rect 300854 57536 300860 57548
rect 300912 57536 300918 57588
rect 320818 57536 320824 57588
rect 320876 57576 320882 57588
rect 444374 57576 444380 57588
rect 320876 57548 444380 57576
rect 320876 57536 320882 57548
rect 444374 57536 444380 57548
rect 444432 57536 444438 57588
rect 449894 57536 449900 57588
rect 449952 57576 449958 57588
rect 450722 57576 450728 57588
rect 449952 57548 450728 57576
rect 449952 57536 449958 57548
rect 450722 57536 450728 57548
rect 450780 57536 450786 57588
rect 452654 57536 452660 57588
rect 452712 57576 452718 57588
rect 453482 57576 453488 57588
rect 452712 57548 453488 57576
rect 452712 57536 452718 57548
rect 453482 57536 453488 57548
rect 453540 57536 453546 57588
rect 455322 57536 455328 57588
rect 455380 57576 455386 57588
rect 484394 57576 484400 57588
rect 455380 57548 484400 57576
rect 455380 57536 455386 57548
rect 484394 57536 484400 57548
rect 484452 57536 484458 57588
rect 497182 57536 497188 57588
rect 497240 57576 497246 57588
rect 498102 57576 498108 57588
rect 497240 57548 498108 57576
rect 497240 57536 497246 57548
rect 498102 57536 498108 57548
rect 498160 57536 498166 57588
rect 516226 57536 516232 57588
rect 516284 57576 516290 57588
rect 517422 57576 517428 57588
rect 516284 57548 517428 57576
rect 516284 57536 516290 57548
rect 517422 57536 517428 57548
rect 517480 57536 517486 57588
rect 140682 57468 140688 57520
rect 140740 57508 140746 57520
rect 171778 57508 171784 57520
rect 140740 57480 171784 57508
rect 140740 57468 140746 57480
rect 171778 57468 171784 57480
rect 171836 57468 171842 57520
rect 183738 57468 183744 57520
rect 183796 57508 183802 57520
rect 184842 57508 184848 57520
rect 183796 57480 184848 57508
rect 183796 57468 183802 57480
rect 184842 57468 184848 57480
rect 184900 57468 184906 57520
rect 186406 57468 186412 57520
rect 186464 57508 186470 57520
rect 187602 57508 187608 57520
rect 186464 57480 187608 57508
rect 186464 57468 186470 57480
rect 187602 57468 187608 57480
rect 187660 57468 187666 57520
rect 190917 57511 190975 57517
rect 190917 57508 190929 57511
rect 190288 57480 190929 57508
rect 133782 57400 133788 57452
rect 133840 57440 133846 57452
rect 170030 57440 170036 57452
rect 133840 57412 170036 57440
rect 133840 57400 133846 57412
rect 170030 57400 170036 57412
rect 170088 57400 170094 57452
rect 188246 57400 188252 57452
rect 188304 57440 188310 57452
rect 190288 57440 190316 57480
rect 190917 57477 190929 57480
rect 190963 57477 190975 57511
rect 190917 57471 190975 57477
rect 191006 57468 191012 57520
rect 191064 57508 191070 57520
rect 191742 57508 191748 57520
rect 191064 57480 191748 57508
rect 191064 57468 191070 57480
rect 191742 57468 191748 57480
rect 191800 57468 191806 57520
rect 191926 57468 191932 57520
rect 191984 57508 191990 57520
rect 193030 57508 193036 57520
rect 191984 57480 193036 57508
rect 191984 57468 191990 57480
rect 193030 57468 193036 57480
rect 193088 57468 193094 57520
rect 193674 57468 193680 57520
rect 193732 57508 193738 57520
rect 194502 57508 194508 57520
rect 193732 57480 194508 57508
rect 193732 57468 193738 57480
rect 194502 57468 194508 57480
rect 194560 57468 194566 57520
rect 194594 57468 194600 57520
rect 194652 57508 194658 57520
rect 195882 57508 195888 57520
rect 194652 57480 195888 57508
rect 194652 57468 194658 57480
rect 195882 57468 195888 57480
rect 195940 57468 195946 57520
rect 196434 57468 196440 57520
rect 196492 57508 196498 57520
rect 197262 57508 197268 57520
rect 196492 57480 197268 57508
rect 196492 57468 196498 57480
rect 197262 57468 197268 57480
rect 197320 57468 197326 57520
rect 197354 57468 197360 57520
rect 197412 57508 197418 57520
rect 198642 57508 198648 57520
rect 197412 57480 198648 57508
rect 197412 57468 197418 57480
rect 198642 57468 198648 57480
rect 198700 57468 198706 57520
rect 199194 57468 199200 57520
rect 199252 57508 199258 57520
rect 200022 57508 200028 57520
rect 199252 57480 200028 57508
rect 199252 57468 199258 57480
rect 200022 57468 200028 57480
rect 200080 57468 200086 57520
rect 200942 57468 200948 57520
rect 201000 57508 201006 57520
rect 201402 57508 201408 57520
rect 201000 57480 201408 57508
rect 201000 57468 201006 57480
rect 201402 57468 201408 57480
rect 201460 57468 201466 57520
rect 201862 57468 201868 57520
rect 201920 57508 201926 57520
rect 202782 57508 202788 57520
rect 201920 57480 202788 57508
rect 201920 57468 201926 57480
rect 202782 57468 202788 57480
rect 202840 57468 202846 57520
rect 203702 57468 203708 57520
rect 203760 57508 203766 57520
rect 204162 57508 204168 57520
rect 203760 57480 204168 57508
rect 203760 57468 203766 57480
rect 204162 57468 204168 57480
rect 204220 57468 204226 57520
rect 204622 57468 204628 57520
rect 204680 57508 204686 57520
rect 205542 57508 205548 57520
rect 204680 57480 205548 57508
rect 204680 57468 204686 57480
rect 205542 57468 205548 57480
rect 205600 57468 205606 57520
rect 206462 57468 206468 57520
rect 206520 57508 206526 57520
rect 206922 57508 206928 57520
rect 206520 57480 206928 57508
rect 206520 57468 206526 57480
rect 206922 57468 206928 57480
rect 206980 57468 206986 57520
rect 209130 57468 209136 57520
rect 209188 57508 209194 57520
rect 209682 57508 209688 57520
rect 209188 57480 209688 57508
rect 209188 57468 209194 57480
rect 209682 57468 209688 57480
rect 209740 57468 209746 57520
rect 212810 57468 212816 57520
rect 212868 57508 212874 57520
rect 213730 57508 213736 57520
rect 212868 57480 213736 57508
rect 212868 57468 212874 57480
rect 213730 57468 213736 57480
rect 213788 57468 213794 57520
rect 214650 57468 214656 57520
rect 214708 57508 214714 57520
rect 215202 57508 215208 57520
rect 214708 57480 215208 57508
rect 214708 57468 214714 57480
rect 215202 57468 215208 57480
rect 215260 57468 215266 57520
rect 215478 57468 215484 57520
rect 215536 57508 215542 57520
rect 216490 57508 216496 57520
rect 215536 57480 216496 57508
rect 215536 57468 215542 57480
rect 216490 57468 216496 57480
rect 216548 57468 216554 57520
rect 217318 57468 217324 57520
rect 217376 57508 217382 57520
rect 217962 57508 217968 57520
rect 217376 57480 217968 57508
rect 217376 57468 217382 57480
rect 217962 57468 217968 57480
rect 218020 57468 218026 57520
rect 219986 57508 219992 57520
rect 218072 57480 219992 57508
rect 188304 57412 190316 57440
rect 190365 57443 190423 57449
rect 188304 57400 188310 57412
rect 190365 57409 190377 57443
rect 190411 57440 190423 57443
rect 200114 57440 200120 57452
rect 190411 57412 200120 57440
rect 190411 57409 190423 57412
rect 190365 57403 190423 57409
rect 200114 57400 200120 57412
rect 200172 57400 200178 57452
rect 211890 57400 211896 57452
rect 211948 57440 211954 57452
rect 218072 57440 218100 57480
rect 219986 57468 219992 57480
rect 220044 57468 220050 57520
rect 220078 57468 220084 57520
rect 220136 57508 220142 57520
rect 220722 57508 220728 57520
rect 220136 57480 220728 57508
rect 220136 57468 220142 57480
rect 220722 57468 220728 57480
rect 220780 57468 220786 57520
rect 222746 57468 222752 57520
rect 222804 57508 222810 57520
rect 223390 57508 223396 57520
rect 222804 57480 223396 57508
rect 222804 57468 222810 57480
rect 223390 57468 223396 57480
rect 223448 57468 223454 57520
rect 223666 57468 223672 57520
rect 223724 57508 223730 57520
rect 224862 57508 224868 57520
rect 223724 57480 224868 57508
rect 223724 57468 223730 57480
rect 224862 57468 224868 57480
rect 224920 57468 224926 57520
rect 229186 57468 229192 57520
rect 229244 57508 229250 57520
rect 230290 57508 230296 57520
rect 229244 57480 230296 57508
rect 229244 57468 229250 57480
rect 230290 57468 230296 57480
rect 230348 57468 230354 57520
rect 230934 57468 230940 57520
rect 230992 57508 230998 57520
rect 231762 57508 231768 57520
rect 230992 57480 231768 57508
rect 230992 57468 230998 57480
rect 231762 57468 231768 57480
rect 231820 57468 231826 57520
rect 231854 57468 231860 57520
rect 231912 57508 231918 57520
rect 233050 57508 233056 57520
rect 231912 57480 233056 57508
rect 231912 57468 231918 57480
rect 233050 57468 233056 57480
rect 233108 57468 233114 57520
rect 233694 57468 233700 57520
rect 233752 57508 233758 57520
rect 234522 57508 234528 57520
rect 233752 57480 234528 57508
rect 233752 57468 233758 57480
rect 234522 57468 234528 57480
rect 234580 57468 234586 57520
rect 237282 57468 237288 57520
rect 237340 57508 237346 57520
rect 238018 57508 238024 57520
rect 237340 57480 238024 57508
rect 237340 57468 237346 57480
rect 238018 57468 238024 57480
rect 238076 57468 238082 57520
rect 384393 57511 384451 57517
rect 384393 57508 384405 57511
rect 238128 57480 384405 57508
rect 211948 57412 218100 57440
rect 211948 57400 211954 57412
rect 219158 57400 219164 57452
rect 219216 57440 219222 57452
rect 221829 57443 221887 57449
rect 221829 57440 221841 57443
rect 219216 57412 221841 57440
rect 219216 57400 219222 57412
rect 221829 57409 221841 57412
rect 221875 57409 221887 57443
rect 221829 57403 221887 57409
rect 221918 57400 221924 57452
rect 221976 57440 221982 57452
rect 231118 57440 231124 57452
rect 221976 57412 231124 57440
rect 221976 57400 221982 57412
rect 231118 57400 231124 57412
rect 231176 57400 231182 57452
rect 236454 57400 236460 57452
rect 236512 57440 236518 57452
rect 238128 57440 238156 57480
rect 384393 57477 384405 57480
rect 384439 57477 384451 57511
rect 384393 57471 384451 57477
rect 384482 57468 384488 57520
rect 384540 57508 384546 57520
rect 384942 57508 384948 57520
rect 384540 57480 384948 57508
rect 384540 57468 384546 57480
rect 384942 57468 384948 57480
rect 385000 57468 385006 57520
rect 385402 57468 385408 57520
rect 385460 57508 385466 57520
rect 386322 57508 386328 57520
rect 385460 57480 386328 57508
rect 385460 57468 385466 57480
rect 386322 57468 386328 57480
rect 386380 57468 386386 57520
rect 387242 57468 387248 57520
rect 387300 57508 387306 57520
rect 387702 57508 387708 57520
rect 387300 57480 387708 57508
rect 387300 57468 387306 57480
rect 387702 57468 387708 57480
rect 387760 57468 387766 57520
rect 388162 57468 388168 57520
rect 388220 57508 388226 57520
rect 388990 57508 388996 57520
rect 388220 57480 388996 57508
rect 388220 57468 388226 57480
rect 388990 57468 388996 57480
rect 389048 57468 389054 57520
rect 390002 57468 390008 57520
rect 390060 57508 390066 57520
rect 390462 57508 390468 57520
rect 390060 57480 390468 57508
rect 390060 57468 390066 57480
rect 390462 57468 390468 57480
rect 390520 57468 390526 57520
rect 390922 57468 390928 57520
rect 390980 57508 390986 57520
rect 391750 57508 391756 57520
rect 390980 57480 391756 57508
rect 390980 57468 390986 57480
rect 391750 57468 391756 57480
rect 391808 57468 391814 57520
rect 392670 57468 392676 57520
rect 392728 57508 392734 57520
rect 393222 57508 393228 57520
rect 392728 57480 393228 57508
rect 392728 57468 392734 57480
rect 393222 57468 393228 57480
rect 393280 57468 393286 57520
rect 393590 57468 393596 57520
rect 393648 57508 393654 57520
rect 394510 57508 394516 57520
rect 393648 57480 394516 57508
rect 393648 57468 393654 57480
rect 394510 57468 394516 57480
rect 394568 57468 394574 57520
rect 395430 57468 395436 57520
rect 395488 57508 395494 57520
rect 395982 57508 395988 57520
rect 395488 57480 395988 57508
rect 395488 57468 395494 57480
rect 395982 57468 395988 57480
rect 396040 57468 396046 57520
rect 396350 57468 396356 57520
rect 396408 57508 396414 57520
rect 397362 57508 397368 57520
rect 396408 57480 397368 57508
rect 396408 57468 396414 57480
rect 397362 57468 397368 57480
rect 397420 57468 397426 57520
rect 398190 57468 398196 57520
rect 398248 57508 398254 57520
rect 398742 57508 398748 57520
rect 398248 57480 398748 57508
rect 398248 57468 398254 57480
rect 398742 57468 398748 57480
rect 398800 57468 398806 57520
rect 399018 57468 399024 57520
rect 399076 57508 399082 57520
rect 400122 57508 400128 57520
rect 399076 57480 400128 57508
rect 399076 57468 399082 57480
rect 400122 57468 400128 57480
rect 400180 57468 400186 57520
rect 404446 57508 404452 57520
rect 402946 57480 404452 57508
rect 236512 57412 238156 57440
rect 236512 57400 236518 57412
rect 238202 57400 238208 57452
rect 238260 57440 238266 57452
rect 238662 57440 238668 57452
rect 238260 57412 238668 57440
rect 238260 57400 238266 57412
rect 238662 57400 238668 57412
rect 238720 57400 238726 57452
rect 240042 57400 240048 57452
rect 240100 57440 240106 57452
rect 240778 57440 240784 57452
rect 240100 57412 240784 57440
rect 240100 57400 240106 57412
rect 240778 57400 240784 57412
rect 240836 57400 240842 57452
rect 240962 57400 240968 57452
rect 241020 57440 241026 57452
rect 241422 57440 241428 57452
rect 241020 57412 241428 57440
rect 241020 57400 241026 57412
rect 241422 57400 241428 57412
rect 241480 57400 241486 57452
rect 241882 57400 241888 57452
rect 241940 57440 241946 57452
rect 242710 57440 242716 57452
rect 241940 57412 242716 57440
rect 241940 57400 241946 57412
rect 242710 57400 242716 57412
rect 242768 57400 242774 57452
rect 243722 57400 243728 57452
rect 243780 57440 243786 57452
rect 244182 57440 244188 57452
rect 243780 57412 244188 57440
rect 243780 57400 243786 57412
rect 244182 57400 244188 57412
rect 244240 57400 244246 57452
rect 244550 57400 244556 57452
rect 244608 57440 244614 57452
rect 245562 57440 245568 57452
rect 244608 57412 245568 57440
rect 244608 57400 244614 57412
rect 245562 57400 245568 57412
rect 245620 57400 245626 57452
rect 246390 57400 246396 57452
rect 246448 57440 246454 57452
rect 246942 57440 246948 57452
rect 246448 57412 246948 57440
rect 246448 57400 246454 57412
rect 246942 57400 246948 57412
rect 247000 57400 247006 57452
rect 247310 57400 247316 57452
rect 247368 57440 247374 57452
rect 248230 57440 248236 57452
rect 247368 57412 248236 57440
rect 247368 57400 247374 57412
rect 248230 57400 248236 57412
rect 248288 57400 248294 57452
rect 248325 57443 248383 57449
rect 248325 57409 248337 57443
rect 248371 57440 248383 57443
rect 394697 57443 394755 57449
rect 394697 57440 394709 57443
rect 248371 57412 394709 57440
rect 248371 57409 248383 57412
rect 248325 57403 248383 57409
rect 394697 57409 394709 57412
rect 394743 57409 394755 57443
rect 394697 57403 394755 57409
rect 394786 57400 394792 57452
rect 394844 57440 394850 57452
rect 402946 57440 402974 57480
rect 404446 57468 404452 57480
rect 404504 57468 404510 57520
rect 412726 57468 412732 57520
rect 412784 57508 412790 57520
rect 413462 57508 413468 57520
rect 412784 57480 413468 57508
rect 412784 57468 412790 57480
rect 413462 57468 413468 57480
rect 413520 57468 413526 57520
rect 415394 57468 415400 57520
rect 415452 57508 415458 57520
rect 416222 57508 416228 57520
rect 415452 57480 416228 57508
rect 415452 57468 415458 57480
rect 416222 57468 416228 57480
rect 416280 57468 416286 57520
rect 418154 57468 418160 57520
rect 418212 57508 418218 57520
rect 418982 57508 418988 57520
rect 418212 57480 418988 57508
rect 418212 57468 418218 57480
rect 418982 57468 418988 57480
rect 419040 57468 419046 57520
rect 435358 57468 435364 57520
rect 435416 57508 435422 57520
rect 440786 57508 440792 57520
rect 435416 57480 440792 57508
rect 435416 57468 435422 57480
rect 440786 57468 440792 57480
rect 440844 57468 440850 57520
rect 448422 57468 448428 57520
rect 448480 57508 448486 57520
rect 482554 57508 482560 57520
rect 448480 57480 482560 57508
rect 448480 57468 448486 57480
rect 482554 57468 482560 57480
rect 482612 57468 482618 57520
rect 394844 57412 402974 57440
rect 394844 57400 394850 57412
rect 403618 57400 403624 57452
rect 403676 57440 403682 57452
rect 438026 57440 438032 57452
rect 403676 57412 438032 57440
rect 403676 57400 403682 57412
rect 438026 57400 438032 57412
rect 438084 57400 438090 57452
rect 441522 57400 441528 57452
rect 441580 57440 441586 57452
rect 480714 57440 480720 57452
rect 441580 57412 480720 57440
rect 441580 57400 441586 57412
rect 480714 57400 480720 57412
rect 480772 57400 480778 57452
rect 487062 57400 487068 57452
rect 487120 57440 487126 57452
rect 492674 57440 492680 57452
rect 487120 57412 492680 57440
rect 487120 57400 487126 57412
rect 492674 57400 492680 57412
rect 492732 57400 492738 57452
rect 501690 57400 501696 57452
rect 501748 57440 501754 57452
rect 502242 57440 502248 57452
rect 501748 57412 502248 57440
rect 501748 57400 501754 57412
rect 502242 57400 502248 57412
rect 502300 57400 502306 57452
rect 504450 57400 504456 57452
rect 504508 57440 504514 57452
rect 505002 57440 505008 57452
rect 504508 57412 505008 57440
rect 504508 57400 504514 57412
rect 505002 57400 505008 57412
rect 505060 57400 505066 57452
rect 507210 57400 507216 57452
rect 507268 57440 507274 57452
rect 507762 57440 507768 57452
rect 507268 57412 507768 57440
rect 507268 57400 507274 57412
rect 507762 57400 507768 57412
rect 507820 57400 507826 57452
rect 2682 57332 2688 57384
rect 2740 57372 2746 57384
rect 72786 57372 72792 57384
rect 2740 57344 72792 57372
rect 2740 57332 2746 57344
rect 72786 57332 72792 57344
rect 72844 57332 72850 57384
rect 129642 57332 129648 57384
rect 129700 57372 129706 57384
rect 169110 57372 169116 57384
rect 129700 57344 169116 57372
rect 129700 57332 129706 57344
rect 169110 57332 169116 57344
rect 169168 57332 169174 57384
rect 188338 57332 188344 57384
rect 188396 57372 188402 57384
rect 408954 57372 408960 57384
rect 188396 57344 408960 57372
rect 188396 57332 188402 57344
rect 408954 57332 408960 57344
rect 409012 57332 409018 57384
rect 421558 57332 421564 57384
rect 421616 57372 421622 57384
rect 427170 57372 427176 57384
rect 421616 57344 427176 57372
rect 421616 57332 421622 57344
rect 427170 57332 427176 57344
rect 427228 57332 427234 57384
rect 433242 57332 433248 57384
rect 433300 57372 433306 57384
rect 478874 57372 478880 57384
rect 433300 57344 478880 57372
rect 433300 57332 433306 57344
rect 478874 57332 478880 57344
rect 478932 57332 478938 57384
rect 480162 57332 480168 57384
rect 480220 57372 480226 57384
rect 490742 57372 490748 57384
rect 480220 57344 490748 57372
rect 480220 57332 480226 57344
rect 490742 57332 490748 57344
rect 490800 57332 490806 57384
rect 491662 57372 491668 57384
rect 490852 57344 491668 57372
rect 126882 57264 126888 57316
rect 126940 57304 126946 57316
rect 168190 57304 168196 57316
rect 126940 57276 168196 57304
rect 126940 57264 126946 57276
rect 168190 57264 168196 57276
rect 168248 57264 168254 57316
rect 173158 57264 173164 57316
rect 173216 57304 173222 57316
rect 407114 57304 407120 57316
rect 173216 57276 407120 57304
rect 173216 57264 173222 57276
rect 407114 57264 407120 57276
rect 407172 57264 407178 57316
rect 423582 57264 423588 57316
rect 423640 57304 423646 57316
rect 476206 57304 476212 57316
rect 423640 57276 476212 57304
rect 423640 57264 423646 57276
rect 476206 57264 476212 57276
rect 476264 57264 476270 57316
rect 482922 57264 482928 57316
rect 482980 57304 482986 57316
rect 490852 57304 490880 57344
rect 491662 57332 491668 57344
rect 491720 57332 491726 57384
rect 482980 57276 490880 57304
rect 482980 57264 482986 57276
rect 491202 57264 491208 57316
rect 491260 57304 491266 57316
rect 493502 57304 493508 57316
rect 491260 57276 493508 57304
rect 491260 57264 491266 57276
rect 493502 57264 493508 57276
rect 493560 57264 493566 57316
rect 1302 57196 1308 57248
rect 1360 57236 1366 57248
rect 72970 57236 72976 57248
rect 1360 57208 72976 57236
rect 1360 57196 1366 57208
rect 72970 57196 72976 57208
rect 73028 57196 73034 57248
rect 162118 57196 162124 57248
rect 162176 57236 162182 57248
rect 405366 57236 405372 57248
rect 162176 57208 405372 57236
rect 162176 57196 162182 57208
rect 405366 57196 405372 57208
rect 405424 57196 405430 57248
rect 416682 57196 416688 57248
rect 416740 57236 416746 57248
rect 474366 57236 474372 57248
rect 416740 57208 474372 57236
rect 416740 57196 416746 57208
rect 474366 57196 474372 57208
rect 474424 57196 474430 57248
rect 476022 57196 476028 57248
rect 476080 57236 476086 57248
rect 489914 57236 489920 57248
rect 476080 57208 489920 57236
rect 476080 57196 476086 57208
rect 489914 57196 489920 57208
rect 489972 57196 489978 57248
rect 169018 57128 169024 57180
rect 169076 57168 169082 57180
rect 287238 57168 287244 57180
rect 169076 57140 287244 57168
rect 169076 57128 169082 57140
rect 287238 57128 287244 57140
rect 287296 57128 287302 57180
rect 382734 57128 382740 57180
rect 382792 57168 382798 57180
rect 383562 57168 383568 57180
rect 382792 57140 383568 57168
rect 382792 57128 382798 57140
rect 383562 57128 383568 57140
rect 383620 57128 383626 57180
rect 384393 57171 384451 57177
rect 384393 57137 384405 57171
rect 384439 57168 384451 57171
rect 389818 57168 389824 57180
rect 384439 57140 389824 57168
rect 384439 57137 384451 57140
rect 384393 57131 384451 57137
rect 389818 57128 389824 57140
rect 389876 57128 389882 57180
rect 394697 57171 394755 57177
rect 394697 57137 394709 57171
rect 394743 57168 394755 57171
rect 400858 57168 400864 57180
rect 394743 57140 400864 57168
rect 394743 57137 394755 57140
rect 394697 57131 394755 57137
rect 400858 57128 400864 57140
rect 400916 57128 400922 57180
rect 144730 57060 144736 57112
rect 144788 57100 144794 57112
rect 172698 57100 172704 57112
rect 144788 57072 172704 57100
rect 144788 57060 144794 57072
rect 172698 57060 172704 57072
rect 172756 57060 172762 57112
rect 189166 57060 189172 57112
rect 189224 57100 189230 57112
rect 190270 57100 190276 57112
rect 189224 57072 190276 57100
rect 189224 57060 189230 57072
rect 190270 57060 190276 57072
rect 190328 57060 190334 57112
rect 190917 57103 190975 57109
rect 190917 57069 190929 57103
rect 190963 57100 190975 57103
rect 196618 57100 196624 57112
rect 190963 57072 196624 57100
rect 190963 57069 190975 57072
rect 190917 57063 190975 57069
rect 196618 57060 196624 57072
rect 196676 57060 196682 57112
rect 210970 57060 210976 57112
rect 211028 57100 211034 57112
rect 211028 57072 258212 57100
rect 211028 57060 211034 57072
rect 151722 56992 151728 57044
rect 151780 57032 151786 57044
rect 174538 57032 174544 57044
rect 151780 57004 174544 57032
rect 151780 56992 151786 57004
rect 174538 56992 174544 57004
rect 174596 56992 174602 57044
rect 207382 56992 207388 57044
rect 207440 57032 207446 57044
rect 208210 57032 208216 57044
rect 207440 57004 208216 57032
rect 207440 56992 207446 57004
rect 208210 56992 208216 57004
rect 208268 56992 208274 57044
rect 210050 56992 210056 57044
rect 210108 57032 210114 57044
rect 214558 57032 214564 57044
rect 210108 57004 214564 57032
rect 210108 56992 210114 57004
rect 214558 56992 214564 57004
rect 214616 56992 214622 57044
rect 221829 57035 221887 57041
rect 221829 57001 221841 57035
rect 221875 57032 221887 57035
rect 228358 57032 228364 57044
rect 221875 57004 228364 57032
rect 221875 57001 221887 57004
rect 221829 56995 221887 57001
rect 228358 56992 228364 57004
rect 228416 56992 228422 57044
rect 239122 56992 239128 57044
rect 239180 57032 239186 57044
rect 248325 57035 248383 57041
rect 248325 57032 248337 57035
rect 239180 57004 248337 57032
rect 239180 56992 239186 57004
rect 248325 57001 248337 57004
rect 248371 57001 248383 57035
rect 248325 56995 248383 57001
rect 249150 56992 249156 57044
rect 249208 57032 249214 57044
rect 249702 57032 249708 57044
rect 249208 57004 249708 57032
rect 249208 56992 249214 57004
rect 249702 56992 249708 57004
rect 249760 56992 249766 57044
rect 250070 56992 250076 57044
rect 250128 57032 250134 57044
rect 250990 57032 250996 57044
rect 250128 57004 250996 57032
rect 250128 56992 250134 57004
rect 250990 56992 250996 57004
rect 251048 56992 251054 57044
rect 251818 56992 251824 57044
rect 251876 57032 251882 57044
rect 252462 57032 252468 57044
rect 251876 57004 252468 57032
rect 251876 56992 251882 57004
rect 252462 56992 252468 57004
rect 252520 56992 252526 57044
rect 252738 56992 252744 57044
rect 252796 57032 252802 57044
rect 253842 57032 253848 57044
rect 252796 57004 253848 57032
rect 252796 56992 252802 57004
rect 253842 56992 253848 57004
rect 253900 56992 253906 57044
rect 254578 56992 254584 57044
rect 254636 57032 254642 57044
rect 255222 57032 255228 57044
rect 254636 57004 255228 57032
rect 254636 56992 254642 57004
rect 255222 56992 255228 57004
rect 255280 56992 255286 57044
rect 255498 56992 255504 57044
rect 255556 57032 255562 57044
rect 256510 57032 256516 57044
rect 255556 57004 256516 57032
rect 255556 56992 255562 57004
rect 256510 56992 256516 57004
rect 256568 56992 256574 57044
rect 257338 56992 257344 57044
rect 257396 57032 257402 57044
rect 257982 57032 257988 57044
rect 257396 57004 257988 57032
rect 257396 56992 257402 57004
rect 257982 56992 257988 57004
rect 258040 56992 258046 57044
rect 258184 57032 258212 57072
rect 258258 57060 258264 57112
rect 258316 57100 258322 57112
rect 259362 57100 259368 57112
rect 258316 57072 259368 57100
rect 258316 57060 258322 57072
rect 259362 57060 259368 57072
rect 259420 57060 259426 57112
rect 260006 57060 260012 57112
rect 260064 57100 260070 57112
rect 260742 57100 260748 57112
rect 260064 57072 260748 57100
rect 260064 57060 260070 57072
rect 260742 57060 260748 57072
rect 260800 57060 260806 57112
rect 262766 57060 262772 57112
rect 262824 57100 262830 57112
rect 263502 57100 263508 57112
rect 262824 57072 263508 57100
rect 262824 57060 262830 57072
rect 263502 57060 263508 57072
rect 263560 57060 263566 57112
rect 263686 57060 263692 57112
rect 263744 57100 263750 57112
rect 264882 57100 264888 57112
rect 263744 57072 264888 57100
rect 263744 57060 263750 57072
rect 264882 57060 264888 57072
rect 264940 57060 264946 57112
rect 266354 57060 266360 57112
rect 266412 57100 266418 57112
rect 267550 57100 267556 57112
rect 266412 57072 267556 57100
rect 266412 57060 266418 57072
rect 267550 57060 267556 57072
rect 267608 57060 267614 57112
rect 268194 57060 268200 57112
rect 268252 57100 268258 57112
rect 269022 57100 269028 57112
rect 268252 57072 269028 57100
rect 268252 57060 268258 57072
rect 269022 57060 269028 57072
rect 269080 57060 269086 57112
rect 269114 57060 269120 57112
rect 269172 57100 269178 57112
rect 270310 57100 270316 57112
rect 269172 57072 270316 57100
rect 269172 57060 269178 57072
rect 270310 57060 270316 57072
rect 270368 57060 270374 57112
rect 270954 57060 270960 57112
rect 271012 57100 271018 57112
rect 271782 57100 271788 57112
rect 271012 57072 271788 57100
rect 271012 57060 271018 57072
rect 271782 57060 271788 57072
rect 271840 57060 271846 57112
rect 271874 57060 271880 57112
rect 271932 57100 271938 57112
rect 273162 57100 273168 57112
rect 271932 57072 273168 57100
rect 271932 57060 271938 57072
rect 273162 57060 273168 57072
rect 273220 57060 273226 57112
rect 273622 57060 273628 57112
rect 273680 57100 273686 57112
rect 274542 57100 274548 57112
rect 273680 57072 274548 57100
rect 273680 57060 273686 57072
rect 274542 57060 274548 57072
rect 274600 57060 274606 57112
rect 275462 57060 275468 57112
rect 275520 57100 275526 57112
rect 275922 57100 275928 57112
rect 275520 57072 275928 57100
rect 275520 57060 275526 57072
rect 275922 57060 275928 57072
rect 275980 57060 275986 57112
rect 276382 57060 276388 57112
rect 276440 57100 276446 57112
rect 277302 57100 277308 57112
rect 276440 57072 277308 57100
rect 276440 57060 276446 57072
rect 277302 57060 277308 57072
rect 277360 57060 277366 57112
rect 278222 57060 278228 57112
rect 278280 57100 278286 57112
rect 278682 57100 278688 57112
rect 278280 57072 278688 57100
rect 278280 57060 278286 57072
rect 278682 57060 278688 57072
rect 278740 57060 278746 57112
rect 279142 57060 279148 57112
rect 279200 57100 279206 57112
rect 279970 57100 279976 57112
rect 279200 57072 279976 57100
rect 279200 57060 279206 57072
rect 279970 57060 279976 57072
rect 280028 57060 280034 57112
rect 280982 57060 280988 57112
rect 281040 57100 281046 57112
rect 281442 57100 281448 57112
rect 281040 57072 281448 57100
rect 281040 57060 281046 57072
rect 281442 57060 281448 57072
rect 281500 57060 281506 57112
rect 281810 57060 281816 57112
rect 281868 57100 281874 57112
rect 282822 57100 282828 57112
rect 281868 57072 282828 57100
rect 281868 57060 281874 57072
rect 282822 57060 282828 57072
rect 282880 57060 282886 57112
rect 283650 57060 283656 57112
rect 283708 57100 283714 57112
rect 284202 57100 284208 57112
rect 283708 57072 284208 57100
rect 283708 57060 283714 57072
rect 284202 57060 284208 57072
rect 284260 57060 284266 57112
rect 286318 57060 286324 57112
rect 286376 57100 286382 57112
rect 319898 57100 319904 57112
rect 286376 57072 319904 57100
rect 286376 57060 286382 57072
rect 319898 57060 319904 57072
rect 319956 57060 319962 57112
rect 264238 57032 264244 57044
rect 258184 57004 264244 57032
rect 264238 56992 264244 57004
rect 264296 56992 264302 57044
rect 287790 57032 287796 57044
rect 264348 57004 287796 57032
rect 147582 56924 147588 56976
rect 147640 56964 147646 56976
rect 173618 56964 173624 56976
rect 147640 56936 173624 56964
rect 147640 56924 147646 56936
rect 173618 56924 173624 56936
rect 173676 56924 173682 56976
rect 259086 56924 259092 56976
rect 259144 56964 259150 56976
rect 264348 56964 264376 57004
rect 287790 56992 287796 57004
rect 287848 56992 287854 57044
rect 288434 56992 288440 57044
rect 288492 57032 288498 57044
rect 292666 57032 292672 57044
rect 288492 57004 292672 57032
rect 288492 56992 288498 57004
rect 292666 56992 292672 57004
rect 292724 56992 292730 57044
rect 259144 56936 264376 56964
rect 259144 56924 259150 56936
rect 264606 56924 264612 56976
rect 264664 56964 264670 56976
rect 291930 56964 291936 56976
rect 264664 56936 291936 56964
rect 264664 56924 264670 56936
rect 291930 56924 291936 56936
rect 291988 56924 291994 56976
rect 158622 56856 158628 56908
rect 158680 56896 158686 56908
rect 176378 56896 176384 56908
rect 158680 56868 176384 56896
rect 158680 56856 158686 56868
rect 176378 56856 176384 56868
rect 176436 56856 176442 56908
rect 228266 56856 228272 56908
rect 228324 56896 228330 56908
rect 229002 56896 229008 56908
rect 228324 56868 229008 56896
rect 228324 56856 228330 56868
rect 229002 56856 229008 56868
rect 229060 56856 229066 56908
rect 289078 56896 289084 56908
rect 277366 56868 289084 56896
rect 161382 56788 161388 56840
rect 161440 56828 161446 56840
rect 177298 56828 177304 56840
rect 161440 56800 177304 56828
rect 161440 56788 161446 56800
rect 177298 56788 177304 56800
rect 177356 56788 177362 56840
rect 165522 56720 165528 56772
rect 165580 56760 165586 56772
rect 178126 56760 178132 56772
rect 165580 56732 178132 56760
rect 165580 56720 165586 56732
rect 178126 56720 178132 56732
rect 178184 56720 178190 56772
rect 260926 56720 260932 56772
rect 260984 56760 260990 56772
rect 277366 56760 277394 56868
rect 289078 56856 289084 56868
rect 289136 56856 289142 56908
rect 260984 56732 277394 56760
rect 260984 56720 260990 56732
rect 309226 56720 309232 56772
rect 309284 56760 309290 56772
rect 309962 56760 309968 56772
rect 309284 56732 309968 56760
rect 309284 56720 309290 56732
rect 309962 56720 309968 56732
rect 310020 56720 310026 56772
rect 347222 56720 347228 56772
rect 347280 56760 347286 56772
rect 347682 56760 347688 56772
rect 347280 56732 347688 56760
rect 347280 56720 347286 56732
rect 347682 56720 347688 56732
rect 347740 56720 347746 56772
rect 349982 56720 349988 56772
rect 350040 56760 350046 56772
rect 350442 56760 350448 56772
rect 350040 56732 350448 56760
rect 350040 56720 350046 56732
rect 350442 56720 350448 56732
rect 350500 56720 350506 56772
rect 352742 56720 352748 56772
rect 352800 56760 352806 56772
rect 353202 56760 353208 56772
rect 352800 56732 353208 56760
rect 352800 56720 352806 56732
rect 353202 56720 353208 56732
rect 353260 56720 353266 56772
rect 361758 56720 361764 56772
rect 361816 56760 361822 56772
rect 362770 56760 362776 56772
rect 361816 56732 362776 56760
rect 361816 56720 361822 56732
rect 362770 56720 362776 56732
rect 362828 56720 362834 56772
rect 166258 56652 166264 56704
rect 166316 56692 166322 56704
rect 175458 56692 175464 56704
rect 166316 56664 175464 56692
rect 166316 56652 166322 56664
rect 175458 56652 175464 56664
rect 175516 56652 175522 56704
rect 178678 56652 178684 56704
rect 178736 56692 178742 56704
rect 180886 56692 180892 56704
rect 178736 56664 180892 56692
rect 178736 56652 178742 56664
rect 180886 56652 180892 56664
rect 180944 56652 180950 56704
rect 185578 56652 185584 56704
rect 185636 56692 185642 56704
rect 191098 56692 191104 56704
rect 185636 56664 191104 56692
rect 185636 56652 185642 56664
rect 191098 56652 191104 56664
rect 191156 56652 191162 56704
rect 180058 56584 180064 56636
rect 180116 56624 180122 56636
rect 181806 56624 181812 56636
rect 180116 56596 181812 56624
rect 180116 56584 180122 56596
rect 181806 56584 181812 56596
rect 181864 56584 181870 56636
rect 220998 56584 221004 56636
rect 221056 56624 221062 56636
rect 221056 56596 223528 56624
rect 221056 56584 221062 56596
rect 223500 56284 223528 56596
rect 287698 56584 287704 56636
rect 287756 56624 287762 56636
rect 288250 56624 288256 56636
rect 287756 56596 288256 56624
rect 287756 56584 287762 56596
rect 288250 56584 288256 56596
rect 288308 56584 288314 56636
rect 291838 56584 291844 56636
rect 291896 56624 291902 56636
rect 297174 56624 297180 56636
rect 291896 56596 297180 56624
rect 291896 56584 291902 56596
rect 297174 56584 297180 56596
rect 297232 56584 297238 56636
rect 429838 56584 429844 56636
rect 429896 56624 429902 56636
rect 434438 56624 434444 56636
rect 429896 56596 434444 56624
rect 429896 56584 429902 56596
rect 434438 56584 434444 56596
rect 434496 56584 434502 56636
rect 262858 56312 262864 56364
rect 262916 56352 262922 56364
rect 318978 56352 318984 56364
rect 262916 56324 318984 56352
rect 262916 56312 262922 56324
rect 318978 56312 318984 56324
rect 319036 56312 319042 56364
rect 382918 56312 382924 56364
rect 382976 56352 382982 56364
rect 456242 56352 456248 56364
rect 382976 56324 456248 56352
rect 382976 56312 382982 56324
rect 456242 56312 456248 56324
rect 456300 56312 456306 56364
rect 331214 56284 331220 56296
rect 223500 56256 331220 56284
rect 331214 56244 331220 56256
rect 331272 56244 331278 56296
rect 363598 56244 363604 56296
rect 363656 56284 363662 56296
rect 451642 56284 451648 56296
rect 363656 56256 451648 56284
rect 363656 56244 363662 56256
rect 451642 56244 451648 56256
rect 451700 56244 451706 56296
rect 177298 56176 177304 56228
rect 177356 56216 177362 56228
rect 294506 56216 294512 56228
rect 177356 56188 294512 56216
rect 177356 56176 177362 56188
rect 294506 56176 294512 56188
rect 294564 56176 294570 56228
rect 322198 56176 322204 56228
rect 322256 56216 322262 56228
rect 441706 56216 441712 56228
rect 322256 56188 441712 56216
rect 322256 56176 322262 56188
rect 441706 56176 441712 56188
rect 441764 56176 441770 56228
rect 170398 56108 170404 56160
rect 170456 56148 170462 56160
rect 293586 56148 293592 56160
rect 170456 56120 293592 56148
rect 170456 56108 170462 56120
rect 293586 56108 293592 56120
rect 293644 56108 293650 56160
rect 318058 56108 318064 56160
rect 318116 56148 318122 56160
rect 445294 56148 445300 56160
rect 318116 56120 445300 56148
rect 318116 56108 318122 56120
rect 445294 56108 445300 56120
rect 445352 56108 445358 56160
rect 447134 56108 447140 56160
rect 447192 56148 447198 56160
rect 448054 56148 448060 56160
rect 447192 56120 448060 56148
rect 447192 56108 447198 56120
rect 448054 56108 448060 56120
rect 448112 56108 448118 56160
rect 280798 56040 280804 56092
rect 280856 56080 280862 56092
rect 433518 56080 433524 56092
rect 280856 56052 433524 56080
rect 280856 56040 280862 56052
rect 433518 56040 433524 56052
rect 433576 56040 433582 56092
rect 261846 55972 261852 56024
rect 261904 56012 261910 56024
rect 489178 56012 489184 56024
rect 261904 55984 489184 56012
rect 261904 55972 261910 55984
rect 489178 55972 489184 55984
rect 489236 55972 489242 56024
rect 265526 55904 265532 55956
rect 265584 55944 265590 55956
rect 504358 55944 504364 55956
rect 265584 55916 504364 55944
rect 265584 55904 265590 55916
rect 504358 55904 504364 55916
rect 504416 55904 504422 55956
rect 137278 55836 137284 55888
rect 137336 55876 137342 55888
rect 402606 55876 402612 55888
rect 137336 55848 402612 55876
rect 137336 55836 137342 55848
rect 402606 55836 402612 55848
rect 402664 55836 402670 55888
rect 298094 55700 298100 55752
rect 298152 55740 298158 55752
rect 299014 55740 299020 55752
rect 298152 55712 299020 55740
rect 298152 55700 298158 55712
rect 299014 55700 299020 55712
rect 299072 55700 299078 55752
rect 226426 54612 226432 54664
rect 226484 54652 226490 54664
rect 351914 54652 351920 54664
rect 226484 54624 351920 54652
rect 226484 54612 226490 54624
rect 351914 54612 351920 54624
rect 351972 54612 351978 54664
rect 160002 54544 160008 54596
rect 160060 54584 160066 54596
rect 288434 54584 288440 54596
rect 160060 54556 288440 54584
rect 160060 54544 160066 54556
rect 288434 54544 288440 54556
rect 288492 54544 288498 54596
rect 340138 54544 340144 54596
rect 340196 54584 340202 54596
rect 447226 54584 447232 54596
rect 340196 54556 447232 54584
rect 340196 54544 340202 54556
rect 447226 54544 447232 54556
rect 447284 54544 447290 54596
rect 143442 54476 143448 54528
rect 143500 54516 143506 54528
rect 394786 54516 394792 54528
rect 143500 54488 394792 54516
rect 143500 54476 143506 54488
rect 394786 54476 394792 54488
rect 394844 54476 394850 54528
rect 233878 50328 233884 50380
rect 233936 50368 233942 50380
rect 349154 50368 349160 50380
rect 233936 50340 349160 50368
rect 233936 50328 233942 50340
rect 349154 50328 349160 50340
rect 349212 50328 349218 50380
rect 522574 46860 522580 46912
rect 522632 46900 522638 46912
rect 580166 46900 580172 46912
rect 522632 46872 580172 46900
rect 522632 46860 522638 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 376018 40672 376024 40724
rect 376076 40712 376082 40724
rect 454034 40712 454040 40724
rect 376076 40684 454040 40712
rect 376076 40672 376082 40684
rect 454034 40672 454040 40684
rect 454092 40672 454098 40724
rect 371878 39312 371884 39364
rect 371936 39352 371942 39364
rect 452746 39352 452752 39364
rect 371936 39324 452752 39352
rect 371936 39312 371942 39324
rect 452746 39312 452752 39324
rect 452804 39312 452810 39364
rect 260098 37884 260104 37936
rect 260156 37924 260162 37936
rect 427906 37924 427912 37936
rect 260156 37896 427912 37924
rect 260156 37884 260162 37896
rect 427906 37884 427912 37896
rect 427964 37884 427970 37936
rect 342898 36524 342904 36576
rect 342956 36564 342962 36576
rect 447134 36564 447140 36576
rect 342956 36536 447140 36564
rect 342956 36524 342962 36536
rect 447134 36524 447140 36536
rect 447192 36524 447198 36576
rect 184198 35164 184204 35216
rect 184256 35204 184262 35216
rect 298186 35204 298192 35216
rect 184256 35176 298192 35204
rect 184256 35164 184262 35176
rect 298186 35164 298192 35176
rect 298244 35164 298250 35216
rect 298738 35164 298744 35216
rect 298796 35204 298802 35216
rect 441614 35204 441620 35216
rect 298796 35176 441620 35204
rect 298796 35164 298802 35176
rect 441614 35164 441620 35176
rect 441672 35164 441678 35216
rect 246298 33736 246304 33788
rect 246356 33776 246362 33788
rect 430666 33776 430672 33788
rect 246356 33748 430672 33776
rect 246356 33736 246362 33748
rect 430666 33736 430672 33748
rect 430724 33736 430730 33788
rect 522482 33056 522488 33108
rect 522540 33096 522546 33108
rect 580166 33096 580172 33108
rect 522540 33068 580172 33096
rect 522540 33056 522546 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 227530 32376 227536 32428
rect 227588 32416 227594 32428
rect 425146 32416 425152 32428
rect 227588 32388 425152 32416
rect 227588 32376 227594 32388
rect 425146 32376 425152 32388
rect 425204 32376 425210 32428
rect 240778 31016 240784 31068
rect 240836 31056 240842 31068
rect 405826 31056 405832 31068
rect 240836 31028 405832 31056
rect 240836 31016 240842 31028
rect 405826 31016 405832 31028
rect 405884 31016 405890 31068
rect 294598 29588 294604 29640
rect 294656 29628 294662 29640
rect 438946 29628 438952 29640
rect 294656 29600 438952 29628
rect 294656 29588 294662 29600
rect 438946 29588 438952 29600
rect 439004 29588 439010 29640
rect 142798 28228 142804 28280
rect 142856 28268 142862 28280
rect 402974 28268 402980 28280
rect 142856 28240 402980 28268
rect 142856 28228 142862 28240
rect 402974 28228 402980 28240
rect 403032 28228 403038 28280
rect 271138 26868 271144 26920
rect 271196 26908 271202 26920
rect 431954 26908 431960 26920
rect 271196 26880 431960 26908
rect 271196 26868 271202 26880
rect 431954 26868 431960 26880
rect 432012 26868 432018 26920
rect 169662 25508 169668 25560
rect 169720 25548 169726 25560
rect 295426 25548 295432 25560
rect 169720 25520 295432 25548
rect 169720 25508 169726 25520
rect 295426 25508 295432 25520
rect 295484 25508 295490 25560
rect 295978 25508 295984 25560
rect 296036 25548 296042 25560
rect 436186 25548 436192 25560
rect 296036 25520 436192 25548
rect 296036 25508 296042 25520
rect 436186 25508 436192 25520
rect 436244 25508 436250 25560
rect 238018 24080 238024 24132
rect 238076 24120 238082 24132
rect 394694 24120 394700 24132
rect 238076 24092 394700 24120
rect 238076 24080 238082 24092
rect 394694 24080 394700 24092
rect 394752 24080 394758 24132
rect 224770 22720 224776 22772
rect 224828 22760 224834 22772
rect 345014 22760 345020 22772
rect 224828 22732 345020 22760
rect 224828 22720 224834 22732
rect 345014 22720 345020 22732
rect 345072 22720 345078 22772
rect 358078 22720 358084 22772
rect 358136 22760 358142 22772
rect 448514 22760 448520 22772
rect 358136 22732 448520 22760
rect 358136 22720 358142 22732
rect 448514 22720 448520 22732
rect 448572 22720 448578 22772
rect 222838 21428 222844 21480
rect 222896 21468 222902 21480
rect 320174 21468 320180 21480
rect 222896 21440 320180 21468
rect 222896 21428 222902 21440
rect 320174 21428 320180 21440
rect 320232 21428 320238 21480
rect 238018 21360 238024 21412
rect 238076 21400 238082 21412
rect 423674 21400 423680 21412
rect 238076 21372 423680 21400
rect 238076 21360 238082 21372
rect 423674 21360 423680 21372
rect 423732 21360 423738 21412
rect 522390 20612 522396 20664
rect 522448 20652 522454 20664
rect 579982 20652 579988 20664
rect 522448 20624 579988 20652
rect 522448 20612 522454 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 268930 20000 268936 20052
rect 268988 20040 268994 20052
rect 320266 20040 320272 20052
rect 268988 20012 320272 20040
rect 268988 20000 268994 20012
rect 320266 20000 320272 20012
rect 320324 20000 320330 20052
rect 214558 19932 214564 19984
rect 214616 19972 214622 19984
rect 288434 19972 288440 19984
rect 214616 19944 288440 19972
rect 214616 19932 214622 19944
rect 288434 19932 288440 19944
rect 288492 19932 288498 19984
rect 323578 19932 323584 19984
rect 323636 19972 323642 19984
rect 442994 19972 443000 19984
rect 323636 19944 443000 19972
rect 323636 19932 323642 19944
rect 442994 19932 443000 19944
rect 443052 19932 443058 19984
rect 357250 18708 357256 18760
rect 357308 18748 357314 18760
rect 407206 18748 407212 18760
rect 357308 18720 407212 18748
rect 357308 18708 357314 18720
rect 407206 18708 407212 18720
rect 407264 18708 407270 18760
rect 231118 18640 231124 18692
rect 231176 18680 231182 18692
rect 334066 18680 334072 18692
rect 231176 18652 334072 18680
rect 231176 18640 231182 18652
rect 334066 18640 334072 18652
rect 334124 18640 334130 18692
rect 356698 18640 356704 18692
rect 356756 18680 356762 18692
rect 449986 18680 449992 18692
rect 356756 18652 449992 18680
rect 356756 18640 356762 18652
rect 449986 18640 449992 18652
rect 450044 18640 450050 18692
rect 231670 18572 231676 18624
rect 231728 18612 231734 18624
rect 421558 18612 421564 18624
rect 231728 18584 421564 18612
rect 231728 18572 231734 18584
rect 421558 18572 421564 18584
rect 421616 18572 421622 18624
rect 214558 17484 214564 17536
rect 214616 17524 214622 17536
rect 299474 17524 299480 17536
rect 214616 17496 299480 17524
rect 214616 17484 214622 17496
rect 299474 17484 299480 17496
rect 299532 17484 299538 17536
rect 378778 17416 378784 17468
rect 378836 17456 378842 17468
rect 456886 17456 456892 17468
rect 378836 17428 456892 17456
rect 378836 17416 378842 17428
rect 456886 17416 456892 17428
rect 456944 17416 456950 17468
rect 213730 17348 213736 17400
rect 213788 17388 213794 17400
rect 299474 17388 299480 17400
rect 213788 17360 299480 17388
rect 213788 17348 213794 17360
rect 299474 17348 299480 17360
rect 299532 17348 299538 17400
rect 379330 17348 379336 17400
rect 379388 17388 379394 17400
rect 486418 17388 486424 17400
rect 379388 17360 486424 17388
rect 379388 17348 379394 17360
rect 486418 17348 486424 17360
rect 486476 17348 486482 17400
rect 298830 17280 298836 17332
rect 298888 17320 298894 17332
rect 434714 17320 434720 17332
rect 298888 17292 434720 17320
rect 298888 17280 298894 17292
rect 434714 17280 434720 17292
rect 434772 17280 434778 17332
rect 278038 17212 278044 17264
rect 278096 17252 278102 17264
rect 436094 17252 436100 17264
rect 278096 17224 436100 17252
rect 278096 17212 278102 17224
rect 436094 17212 436100 17224
rect 436152 17212 436158 17264
rect 224218 16124 224224 16176
rect 224276 16164 224282 16176
rect 298094 16164 298100 16176
rect 224276 16136 298100 16164
rect 224276 16124 224282 16136
rect 298094 16124 298100 16136
rect 298152 16124 298158 16176
rect 266998 16056 267004 16108
rect 267056 16096 267062 16108
rect 430574 16096 430580 16108
rect 267056 16068 430580 16096
rect 267056 16056 267062 16068
rect 430574 16056 430580 16068
rect 430632 16056 430638 16108
rect 249058 15988 249064 16040
rect 249116 16028 249122 16040
rect 427814 16028 427820 16040
rect 249116 16000 427820 16028
rect 249116 15988 249122 16000
rect 427814 15988 427820 16000
rect 427872 15988 427878 16040
rect 228450 15920 228456 15972
rect 228508 15960 228514 15972
rect 425054 15960 425060 15972
rect 228508 15932 425060 15960
rect 228508 15920 228514 15932
rect 425054 15920 425060 15932
rect 425112 15920 425118 15972
rect 267550 15852 267556 15904
rect 267608 15892 267614 15904
rect 507118 15892 507124 15904
rect 267608 15864 507124 15892
rect 267608 15852 267614 15864
rect 507118 15852 507124 15864
rect 507176 15852 507182 15904
rect 259270 14900 259276 14952
rect 259328 14940 259334 14952
rect 317414 14940 317420 14952
rect 259328 14912 317420 14940
rect 259328 14900 259334 14912
rect 317414 14900 317420 14912
rect 317472 14900 317478 14952
rect 173802 14832 173808 14884
rect 173860 14872 173866 14884
rect 295334 14872 295340 14884
rect 173860 14844 295340 14872
rect 173860 14832 173866 14844
rect 295334 14832 295340 14844
rect 295392 14832 295398 14884
rect 318150 14832 318156 14884
rect 318208 14872 318214 14884
rect 438854 14872 438860 14884
rect 318208 14844 438860 14872
rect 318208 14832 318214 14844
rect 438854 14832 438860 14844
rect 438912 14832 438918 14884
rect 274358 14764 274364 14816
rect 274416 14804 274422 14816
rect 403618 14804 403624 14816
rect 274416 14776 403624 14804
rect 274416 14764 274422 14776
rect 403618 14764 403624 14776
rect 403676 14764 403682 14816
rect 229002 14696 229008 14748
rect 229060 14736 229066 14748
rect 359458 14736 359464 14748
rect 229060 14708 359464 14736
rect 229060 14696 229066 14708
rect 359458 14696 359464 14708
rect 359516 14696 359522 14748
rect 360838 14696 360844 14748
rect 360896 14736 360902 14748
rect 449894 14736 449900 14748
rect 360896 14708 449900 14736
rect 360896 14696 360902 14708
rect 449894 14696 449900 14708
rect 449952 14696 449958 14748
rect 242710 14628 242716 14680
rect 242768 14668 242774 14680
rect 412634 14668 412640 14680
rect 242768 14640 412640 14668
rect 242768 14628 242774 14640
rect 412634 14628 412640 14640
rect 412692 14628 412698 14680
rect 235902 14560 235908 14612
rect 235960 14600 235966 14612
rect 387794 14600 387800 14612
rect 235960 14572 387800 14600
rect 235960 14560 235966 14572
rect 387794 14560 387800 14572
rect 387852 14560 387858 14612
rect 242710 14492 242716 14544
rect 242768 14532 242774 14544
rect 429194 14532 429200 14544
rect 242768 14504 429200 14532
rect 242768 14492 242774 14504
rect 429194 14492 429200 14504
rect 429252 14492 429258 14544
rect 264882 14424 264888 14476
rect 264940 14464 264946 14476
rect 490558 14464 490564 14476
rect 264940 14436 490564 14464
rect 264940 14424 264946 14436
rect 490558 14424 490564 14436
rect 490616 14424 490622 14476
rect 255958 13676 255964 13728
rect 256016 13716 256022 13728
rect 316126 13716 316132 13728
rect 256016 13688 316132 13716
rect 256016 13676 256022 13688
rect 316126 13676 316132 13688
rect 316184 13676 316190 13728
rect 228358 13608 228364 13660
rect 228416 13648 228422 13660
rect 324406 13648 324412 13660
rect 228416 13620 324412 13648
rect 228416 13608 228422 13620
rect 324406 13608 324412 13620
rect 324464 13608 324470 13660
rect 217962 13540 217968 13592
rect 218020 13580 218026 13592
rect 317322 13580 317328 13592
rect 218020 13552 317328 13580
rect 218020 13540 218026 13552
rect 317322 13540 317328 13552
rect 317380 13540 317386 13592
rect 383562 13540 383568 13592
rect 383620 13580 383626 13592
rect 467098 13580 467104 13592
rect 383620 13552 467104 13580
rect 383620 13540 383626 13552
rect 467098 13540 467104 13552
rect 467156 13540 467162 13592
rect 224862 13472 224868 13524
rect 224920 13512 224926 13524
rect 340874 13512 340880 13524
rect 224920 13484 340880 13512
rect 224920 13472 224926 13484
rect 340874 13472 340880 13484
rect 340932 13472 340938 13524
rect 378042 13472 378048 13524
rect 378100 13512 378106 13524
rect 488810 13512 488816 13524
rect 378100 13484 488816 13512
rect 378100 13472 378106 13484
rect 488810 13472 488816 13484
rect 488868 13472 488874 13524
rect 220722 13404 220728 13456
rect 220780 13444 220786 13456
rect 327074 13444 327080 13456
rect 220780 13416 327080 13444
rect 220780 13404 220786 13416
rect 327074 13404 327080 13416
rect 327132 13404 327138 13456
rect 334710 13404 334716 13456
rect 334768 13444 334774 13456
rect 452654 13444 452660 13456
rect 334768 13416 452660 13444
rect 334768 13404 334774 13416
rect 452654 13404 452660 13416
rect 452712 13404 452718 13456
rect 285582 13336 285588 13388
rect 285640 13376 285646 13388
rect 435358 13376 435364 13388
rect 285640 13348 435364 13376
rect 285640 13336 285646 13348
rect 435358 13336 435364 13348
rect 435416 13336 435422 13388
rect 238662 13268 238668 13320
rect 238720 13308 238726 13320
rect 398926 13308 398932 13320
rect 238720 13280 398932 13308
rect 238720 13268 238726 13280
rect 398926 13268 398932 13280
rect 398984 13268 398990 13320
rect 260650 13200 260656 13252
rect 260708 13240 260714 13252
rect 429838 13240 429844 13252
rect 260708 13212 429844 13240
rect 260708 13200 260714 13212
rect 429838 13200 429844 13212
rect 429896 13200 429902 13252
rect 291930 13132 291936 13184
rect 291988 13172 291994 13184
rect 501322 13172 501328 13184
rect 291988 13144 501328 13172
rect 291988 13132 291994 13144
rect 501322 13132 501328 13144
rect 501380 13132 501386 13184
rect 263502 13064 263508 13116
rect 263560 13104 263566 13116
rect 493318 13104 493324 13116
rect 263560 13076 493324 13104
rect 263560 13064 263566 13076
rect 493318 13064 493324 13076
rect 493376 13064 493382 13116
rect 277118 12384 277124 12436
rect 277176 12424 277182 12436
rect 321646 12424 321652 12436
rect 277176 12396 321652 12424
rect 277176 12384 277182 12396
rect 321646 12384 321652 12396
rect 321704 12384 321710 12436
rect 215202 12316 215208 12368
rect 215260 12356 215266 12368
rect 306374 12356 306380 12368
rect 215260 12328 306380 12356
rect 215260 12316 215266 12328
rect 306374 12316 306380 12328
rect 306432 12316 306438 12368
rect 216490 12248 216496 12300
rect 216548 12288 216554 12300
rect 309778 12288 309784 12300
rect 216548 12260 309784 12288
rect 216548 12248 216554 12260
rect 309778 12248 309784 12260
rect 309836 12248 309842 12300
rect 357342 12248 357348 12300
rect 357400 12288 357406 12300
rect 410794 12288 410800 12300
rect 357400 12260 410800 12288
rect 357400 12248 357406 12260
rect 410794 12248 410800 12260
rect 410852 12248 410858 12300
rect 216582 12180 216588 12232
rect 216640 12220 216646 12232
rect 313826 12220 313832 12232
rect 216640 12192 313832 12220
rect 216640 12180 216646 12192
rect 313826 12180 313832 12192
rect 313884 12180 313890 12232
rect 376662 12180 376668 12232
rect 376720 12220 376726 12232
rect 484486 12220 484492 12232
rect 376720 12192 484492 12220
rect 376720 12180 376726 12192
rect 484486 12180 484492 12192
rect 484544 12180 484550 12232
rect 223482 12112 223488 12164
rect 223540 12152 223546 12164
rect 338666 12152 338672 12164
rect 223540 12124 338672 12152
rect 223540 12112 223546 12124
rect 338666 12112 338672 12124
rect 338724 12112 338730 12164
rect 379422 12112 379428 12164
rect 379480 12152 379486 12164
rect 495434 12152 495440 12164
rect 379480 12124 495440 12152
rect 379480 12112 379486 12124
rect 495434 12112 495440 12124
rect 495492 12112 495498 12164
rect 227622 12044 227628 12096
rect 227680 12084 227686 12096
rect 356330 12084 356336 12096
rect 227680 12056 356336 12084
rect 227680 12044 227686 12056
rect 356330 12044 356336 12056
rect 356388 12044 356394 12096
rect 382182 12044 382188 12096
rect 382240 12084 382246 12096
rect 506474 12084 506480 12096
rect 382240 12056 506480 12084
rect 382240 12044 382246 12056
rect 506474 12044 506480 12056
rect 506532 12044 506538 12096
rect 213822 11976 213828 12028
rect 213880 12016 213886 12028
rect 303154 12016 303160 12028
rect 213880 11988 303160 12016
rect 213880 11976 213886 11988
rect 303154 11976 303160 11988
rect 303212 11976 303218 12028
rect 306282 11976 306288 12028
rect 306340 12016 306346 12028
rect 445754 12016 445760 12028
rect 306340 11988 445760 12016
rect 306340 11976 306346 11988
rect 445754 11976 445760 11988
rect 445812 11976 445818 12028
rect 241422 11908 241428 11960
rect 241480 11948 241486 11960
rect 409138 11948 409144 11960
rect 241480 11920 409144 11948
rect 241480 11908 241486 11920
rect 409138 11908 409144 11920
rect 409196 11908 409202 11960
rect 287790 11840 287796 11892
rect 287848 11880 287854 11892
rect 480530 11880 480536 11892
rect 287848 11852 480536 11880
rect 287848 11840 287854 11852
rect 480530 11840 480536 11852
rect 480588 11840 480594 11892
rect 289078 11772 289084 11824
rect 289136 11812 289142 11824
rect 487154 11812 487160 11824
rect 289136 11784 487160 11812
rect 289136 11772 289142 11784
rect 487154 11772 487160 11784
rect 487212 11772 487218 11824
rect 260742 11704 260748 11756
rect 260800 11744 260806 11756
rect 483658 11744 483664 11756
rect 260800 11716 483664 11744
rect 260800 11704 260806 11716
rect 483658 11704 483664 11716
rect 483716 11704 483722 11756
rect 192938 10956 192944 11008
rect 192996 10996 193002 11008
rect 416774 10996 416780 11008
rect 192996 10968 416780 10996
rect 192996 10956 193002 10968
rect 416774 10956 416780 10968
rect 416832 10956 416838 11008
rect 188982 10888 188988 10940
rect 189040 10928 189046 10940
rect 415394 10928 415400 10940
rect 189040 10900 415400 10928
rect 189040 10888 189046 10900
rect 415394 10888 415400 10900
rect 415452 10888 415458 10940
rect 186222 10820 186228 10872
rect 186280 10860 186286 10872
rect 415486 10860 415492 10872
rect 186280 10832 415492 10860
rect 186280 10820 186286 10832
rect 415486 10820 415492 10832
rect 415544 10820 415550 10872
rect 182082 10752 182088 10804
rect 182140 10792 182146 10804
rect 414014 10792 414020 10804
rect 182140 10764 414020 10792
rect 182140 10752 182146 10764
rect 414014 10752 414020 10764
rect 414072 10752 414078 10804
rect 177850 10684 177856 10736
rect 177908 10724 177914 10736
rect 412726 10724 412732 10736
rect 177908 10696 412732 10724
rect 177908 10684 177914 10696
rect 412726 10684 412732 10696
rect 412784 10684 412790 10736
rect 175182 10616 175188 10668
rect 175240 10656 175246 10668
rect 412818 10656 412824 10668
rect 175240 10628 412824 10656
rect 175240 10616 175246 10628
rect 412818 10616 412824 10628
rect 412876 10616 412882 10668
rect 170766 10548 170772 10600
rect 170824 10588 170830 10600
rect 411254 10588 411260 10600
rect 170824 10560 411260 10588
rect 170824 10548 170830 10560
rect 411254 10548 411260 10560
rect 411312 10548 411318 10600
rect 168282 10480 168288 10532
rect 168340 10520 168346 10532
rect 410058 10520 410064 10532
rect 168340 10492 410064 10520
rect 168340 10480 168346 10492
rect 410058 10480 410064 10492
rect 410116 10480 410122 10532
rect 164142 10412 164148 10464
rect 164200 10452 164206 10464
rect 409966 10452 409972 10464
rect 164200 10424 409972 10452
rect 164200 10412 164206 10424
rect 409966 10412 409972 10424
rect 410024 10412 410030 10464
rect 132402 10344 132408 10396
rect 132460 10384 132466 10396
rect 401594 10384 401600 10396
rect 132460 10356 401600 10384
rect 132460 10344 132466 10356
rect 401594 10344 401600 10356
rect 401652 10344 401658 10396
rect 128170 10276 128176 10328
rect 128228 10316 128234 10328
rect 400214 10316 400220 10328
rect 128228 10288 400220 10316
rect 128228 10276 128234 10288
rect 400214 10276 400220 10288
rect 400272 10276 400278 10328
rect 195606 10208 195612 10260
rect 195664 10248 195670 10260
rect 418246 10248 418252 10260
rect 195664 10220 418252 10248
rect 195664 10208 195670 10220
rect 418246 10208 418252 10220
rect 418304 10208 418310 10260
rect 199930 10140 199936 10192
rect 199988 10180 199994 10192
rect 418154 10180 418160 10192
rect 199988 10152 418160 10180
rect 199988 10140 199994 10152
rect 418154 10140 418160 10152
rect 418212 10140 418218 10192
rect 202598 10072 202604 10124
rect 202656 10112 202662 10124
rect 419534 10112 419540 10124
rect 202656 10084 419540 10112
rect 202656 10072 202662 10084
rect 419534 10072 419540 10084
rect 419592 10072 419598 10124
rect 206830 10004 206836 10056
rect 206888 10044 206894 10056
rect 419626 10044 419632 10056
rect 206888 10016 419632 10044
rect 206888 10004 206894 10016
rect 419626 10004 419632 10016
rect 419684 10004 419690 10056
rect 211062 9936 211068 9988
rect 211120 9976 211126 9988
rect 420914 9976 420920 9988
rect 211120 9948 420920 9976
rect 211120 9936 211126 9948
rect 420914 9936 420920 9948
rect 420972 9936 420978 9988
rect 213822 9868 213828 9920
rect 213880 9908 213886 9920
rect 422294 9908 422300 9920
rect 213880 9880 422300 9908
rect 213880 9868 213886 9880
rect 422294 9868 422300 9880
rect 422352 9868 422358 9920
rect 217962 9800 217968 9852
rect 218020 9840 218026 9852
rect 422386 9840 422392 9852
rect 218020 9812 422392 9840
rect 218020 9800 218026 9812
rect 422386 9800 422392 9812
rect 422444 9800 422450 9852
rect 284110 9732 284116 9784
rect 284168 9772 284174 9784
rect 324498 9772 324504 9784
rect 284168 9744 324504 9772
rect 284168 9732 284174 9744
rect 324498 9732 324504 9744
rect 324556 9732 324562 9784
rect 222746 9596 222752 9648
rect 222804 9636 222810 9648
rect 309318 9636 309324 9648
rect 222804 9608 309324 9636
rect 222804 9596 222810 9608
rect 309318 9596 309324 9608
rect 309376 9596 309382 9648
rect 365622 9596 365628 9648
rect 365680 9636 365686 9648
rect 442626 9636 442632 9648
rect 365680 9608 442632 9636
rect 365680 9596 365686 9608
rect 442626 9596 442632 9608
rect 442684 9596 442690 9648
rect 449802 9636 449808 9648
rect 446324 9608 449808 9636
rect 219250 9528 219256 9580
rect 219308 9568 219314 9580
rect 307754 9568 307760 9580
rect 219308 9540 307760 9568
rect 219308 9528 219314 9540
rect 307754 9528 307760 9540
rect 307812 9528 307818 9580
rect 367002 9528 367008 9580
rect 367060 9568 367066 9580
rect 446214 9568 446220 9580
rect 367060 9540 446220 9568
rect 367060 9528 367066 9540
rect 446214 9528 446220 9540
rect 446272 9528 446278 9580
rect 215662 9460 215668 9512
rect 215720 9500 215726 9512
rect 306558 9500 306564 9512
rect 215720 9472 306564 9500
rect 215720 9460 215726 9472
rect 306558 9460 306564 9472
rect 306616 9460 306622 9512
rect 368382 9460 368388 9512
rect 368440 9500 368446 9512
rect 446324 9500 446352 9608
rect 449802 9596 449808 9608
rect 449860 9596 449866 9648
rect 453298 9568 453304 9580
rect 368440 9472 446352 9500
rect 446416 9540 453304 9568
rect 368440 9460 368446 9472
rect 212166 9392 212172 9444
rect 212224 9432 212230 9444
rect 306466 9432 306472 9444
rect 212224 9404 306472 9432
rect 212224 9392 212230 9404
rect 306466 9392 306472 9404
rect 306524 9392 306530 9444
rect 368290 9392 368296 9444
rect 368348 9432 368354 9444
rect 446416 9432 446444 9540
rect 453298 9528 453304 9540
rect 453356 9528 453362 9580
rect 449158 9460 449164 9512
rect 449216 9500 449222 9512
rect 502978 9500 502984 9512
rect 449216 9472 502984 9500
rect 449216 9460 449222 9472
rect 502978 9460 502984 9472
rect 503036 9460 503042 9512
rect 368348 9404 446444 9432
rect 368348 9392 368354 9404
rect 208578 9324 208584 9376
rect 208636 9364 208642 9376
rect 304994 9364 305000 9376
rect 208636 9336 305000 9364
rect 208636 9324 208642 9336
rect 304994 9324 305000 9336
rect 305052 9324 305058 9376
rect 369762 9324 369768 9376
rect 369820 9364 369826 9376
rect 456886 9364 456892 9376
rect 369820 9336 456892 9364
rect 369820 9324 369826 9336
rect 456886 9324 456892 9336
rect 456944 9324 456950 9376
rect 205082 9256 205088 9308
rect 205140 9296 205146 9308
rect 303706 9296 303712 9308
rect 205140 9268 303712 9296
rect 205140 9256 205146 9268
rect 303706 9256 303712 9268
rect 303764 9256 303770 9308
rect 371050 9256 371056 9308
rect 371108 9296 371114 9308
rect 460382 9296 460388 9308
rect 371108 9268 460388 9296
rect 371108 9256 371114 9268
rect 460382 9256 460388 9268
rect 460440 9256 460446 9308
rect 201494 9188 201500 9240
rect 201552 9228 201558 9240
rect 303614 9228 303620 9240
rect 201552 9200 303620 9228
rect 201552 9188 201558 9200
rect 303614 9188 303620 9200
rect 303672 9188 303678 9240
rect 371142 9188 371148 9240
rect 371200 9228 371206 9240
rect 463970 9228 463976 9240
rect 371200 9200 463976 9228
rect 371200 9188 371206 9200
rect 463970 9188 463976 9200
rect 464028 9188 464034 9240
rect 197906 9120 197912 9172
rect 197964 9160 197970 9172
rect 302326 9160 302332 9172
rect 197964 9132 302332 9160
rect 197964 9120 197970 9132
rect 302326 9120 302332 9132
rect 302384 9120 302390 9172
rect 372522 9120 372528 9172
rect 372580 9160 372586 9172
rect 467466 9160 467472 9172
rect 372580 9132 467472 9160
rect 372580 9120 372586 9132
rect 467466 9120 467472 9132
rect 467524 9120 467530 9172
rect 194410 9052 194416 9104
rect 194468 9092 194474 9104
rect 300946 9092 300952 9104
rect 194468 9064 300952 9092
rect 194468 9052 194474 9064
rect 300946 9052 300952 9064
rect 301004 9052 301010 9104
rect 373810 9052 373816 9104
rect 373868 9092 373874 9104
rect 471054 9092 471060 9104
rect 373868 9064 471060 9092
rect 373868 9052 373874 9064
rect 471054 9052 471060 9064
rect 471112 9052 471118 9104
rect 134150 8984 134156 9036
rect 134208 9024 134214 9036
rect 285674 9024 285680 9036
rect 134208 8996 285680 9024
rect 134208 8984 134214 8996
rect 285674 8984 285680 8996
rect 285732 8984 285738 9036
rect 373902 8984 373908 9036
rect 373960 9024 373966 9036
rect 474550 9024 474556 9036
rect 373960 8996 474556 9024
rect 373960 8984 373966 8996
rect 474550 8984 474556 8996
rect 474608 8984 474614 9036
rect 130562 8916 130568 8968
rect 130620 8956 130626 8968
rect 284386 8956 284392 8968
rect 130620 8928 284392 8956
rect 130620 8916 130626 8928
rect 284386 8916 284392 8928
rect 284444 8916 284450 8968
rect 375282 8916 375288 8968
rect 375340 8956 375346 8968
rect 478138 8956 478144 8968
rect 375340 8928 478144 8956
rect 375340 8916 375346 8928
rect 478138 8916 478144 8928
rect 478196 8916 478202 8968
rect 226334 8848 226340 8900
rect 226392 8888 226398 8900
rect 309226 8888 309232 8900
rect 226392 8860 309232 8888
rect 226392 8848 226398 8860
rect 309226 8848 309232 8860
rect 309284 8848 309290 8900
rect 365530 8848 365536 8900
rect 365588 8888 365594 8900
rect 439130 8888 439136 8900
rect 365588 8860 439136 8888
rect 365588 8848 365594 8860
rect 439130 8848 439136 8860
rect 439188 8848 439194 8900
rect 229830 8780 229836 8832
rect 229888 8820 229894 8832
rect 310514 8820 310520 8832
rect 229888 8792 310520 8820
rect 229888 8780 229894 8792
rect 310514 8780 310520 8792
rect 310572 8780 310578 8832
rect 364242 8780 364248 8832
rect 364300 8820 364306 8832
rect 435542 8820 435548 8832
rect 364300 8792 435548 8820
rect 364300 8780 364306 8792
rect 435542 8780 435548 8792
rect 435600 8780 435606 8832
rect 233418 8712 233424 8764
rect 233476 8752 233482 8764
rect 310606 8752 310612 8764
rect 233476 8724 310612 8752
rect 233476 8712 233482 8724
rect 310606 8712 310612 8724
rect 310664 8712 310670 8764
rect 362862 8712 362868 8764
rect 362920 8752 362926 8764
rect 432046 8752 432052 8764
rect 362920 8724 432052 8752
rect 362920 8712 362926 8724
rect 432046 8712 432052 8724
rect 432104 8712 432110 8764
rect 237006 8644 237012 8696
rect 237064 8684 237070 8696
rect 311894 8684 311900 8696
rect 237064 8656 311900 8684
rect 237064 8644 237070 8656
rect 311894 8644 311900 8656
rect 311952 8644 311958 8696
rect 362770 8644 362776 8696
rect 362828 8684 362834 8696
rect 428458 8684 428464 8696
rect 362828 8656 428464 8684
rect 362828 8644 362834 8656
rect 428458 8644 428464 8656
rect 428516 8644 428522 8696
rect 240502 8576 240508 8628
rect 240560 8616 240566 8628
rect 313458 8616 313464 8628
rect 240560 8588 313464 8616
rect 240560 8576 240566 8588
rect 313458 8576 313464 8588
rect 313516 8576 313522 8628
rect 361482 8576 361488 8628
rect 361540 8616 361546 8628
rect 424962 8616 424968 8628
rect 361540 8588 424968 8616
rect 361540 8576 361546 8588
rect 424962 8576 424968 8588
rect 425020 8576 425026 8628
rect 244090 8508 244096 8560
rect 244148 8548 244154 8560
rect 313366 8548 313372 8560
rect 244148 8520 313372 8548
rect 244148 8508 244154 8520
rect 313366 8508 313372 8520
rect 313424 8508 313430 8560
rect 360102 8508 360108 8560
rect 360160 8548 360166 8560
rect 421374 8548 421380 8560
rect 360160 8520 421380 8548
rect 360160 8508 360166 8520
rect 421374 8508 421380 8520
rect 421432 8508 421438 8560
rect 247586 8440 247592 8492
rect 247644 8480 247650 8492
rect 314654 8480 314660 8492
rect 247644 8452 314660 8480
rect 247644 8440 247650 8452
rect 314654 8440 314660 8452
rect 314712 8440 314718 8492
rect 360010 8440 360016 8492
rect 360068 8480 360074 8492
rect 417878 8480 417884 8492
rect 360068 8452 417884 8480
rect 360068 8440 360074 8452
rect 417878 8440 417884 8452
rect 417936 8440 417942 8492
rect 251174 8372 251180 8424
rect 251232 8412 251238 8424
rect 316034 8412 316040 8424
rect 251232 8384 316040 8412
rect 251232 8372 251238 8384
rect 316034 8372 316040 8384
rect 316092 8372 316098 8424
rect 358722 8372 358728 8424
rect 358780 8412 358786 8424
rect 414290 8412 414296 8424
rect 358780 8384 414296 8412
rect 358780 8372 358786 8384
rect 414290 8372 414296 8384
rect 414348 8372 414354 8424
rect 249702 8236 249708 8288
rect 249760 8276 249766 8288
rect 441246 8276 441252 8288
rect 249760 8248 441252 8276
rect 249760 8236 249766 8248
rect 441246 8236 441252 8248
rect 441304 8236 441310 8288
rect 443638 8236 443644 8288
rect 443696 8276 443702 8288
rect 481726 8276 481732 8288
rect 443696 8248 481732 8276
rect 443696 8236 443702 8248
rect 481726 8236 481732 8248
rect 481784 8236 481790 8288
rect 250990 8168 250996 8220
rect 251048 8208 251054 8220
rect 445018 8208 445024 8220
rect 251048 8180 445024 8208
rect 251048 8168 251054 8180
rect 445018 8168 445024 8180
rect 445076 8168 445082 8220
rect 251082 8100 251088 8152
rect 251140 8140 251146 8152
rect 448606 8140 448612 8152
rect 251140 8112 448612 8140
rect 251140 8100 251146 8112
rect 448606 8100 448612 8112
rect 448664 8100 448670 8152
rect 252462 8032 252468 8084
rect 252520 8072 252526 8084
rect 452102 8072 452108 8084
rect 252520 8044 452108 8072
rect 252520 8032 252526 8044
rect 452102 8032 452108 8044
rect 452160 8032 452166 8084
rect 253842 7964 253848 8016
rect 253900 8004 253906 8016
rect 455690 8004 455696 8016
rect 253900 7976 455696 8004
rect 253900 7964 253906 7976
rect 455690 7964 455696 7976
rect 455748 7964 455754 8016
rect 253750 7896 253756 7948
rect 253808 7936 253814 7948
rect 459186 7936 459192 7948
rect 253808 7908 459192 7936
rect 253808 7896 253814 7908
rect 459186 7896 459192 7908
rect 459244 7896 459250 7948
rect 255222 7828 255228 7880
rect 255280 7868 255286 7880
rect 462774 7868 462780 7880
rect 255280 7840 462780 7868
rect 255280 7828 255286 7840
rect 462774 7828 462780 7840
rect 462832 7828 462838 7880
rect 256510 7760 256516 7812
rect 256568 7800 256574 7812
rect 466270 7800 466276 7812
rect 256568 7772 466276 7800
rect 256568 7760 256574 7772
rect 466270 7760 466276 7772
rect 466328 7760 466334 7812
rect 256602 7692 256608 7744
rect 256660 7732 256666 7744
rect 469858 7732 469864 7744
rect 256660 7704 469864 7732
rect 256660 7692 256666 7704
rect 469858 7692 469864 7704
rect 469916 7692 469922 7744
rect 257982 7624 257988 7676
rect 258040 7664 258046 7676
rect 473446 7664 473452 7676
rect 258040 7636 473452 7664
rect 258040 7624 258046 7636
rect 473446 7624 473452 7636
rect 473504 7624 473510 7676
rect 259362 7556 259368 7608
rect 259420 7596 259426 7608
rect 476942 7596 476948 7608
rect 259420 7568 476948 7596
rect 259420 7556 259426 7568
rect 476942 7556 476948 7568
rect 477000 7556 477006 7608
rect 248322 7488 248328 7540
rect 248380 7528 248386 7540
rect 437934 7528 437940 7540
rect 248380 7500 437940 7528
rect 248380 7488 248386 7500
rect 437934 7488 437940 7500
rect 437992 7488 437998 7540
rect 248230 7420 248236 7472
rect 248288 7460 248294 7472
rect 434438 7460 434444 7472
rect 248288 7432 434444 7460
rect 248288 7420 248294 7432
rect 434438 7420 434444 7432
rect 434496 7420 434502 7472
rect 246942 7352 246948 7404
rect 247000 7392 247006 7404
rect 430850 7392 430856 7404
rect 247000 7364 430856 7392
rect 247000 7352 247006 7364
rect 430850 7352 430856 7364
rect 430908 7352 430914 7404
rect 245470 7284 245476 7336
rect 245528 7324 245534 7336
rect 427262 7324 427268 7336
rect 245528 7296 427268 7324
rect 245528 7284 245534 7296
rect 427262 7284 427268 7296
rect 427320 7284 427326 7336
rect 245562 7216 245568 7268
rect 245620 7256 245626 7268
rect 423766 7256 423772 7268
rect 245620 7228 423772 7256
rect 245620 7216 245626 7228
rect 423766 7216 423772 7228
rect 423824 7216 423830 7268
rect 244182 7148 244188 7200
rect 244240 7188 244246 7200
rect 420178 7188 420184 7200
rect 244240 7160 420184 7188
rect 244240 7148 244246 7160
rect 420178 7148 420184 7160
rect 420236 7148 420242 7200
rect 242802 7080 242808 7132
rect 242860 7120 242866 7132
rect 416406 7120 416412 7132
rect 242860 7092 416412 7120
rect 242860 7080 242866 7092
rect 416406 7080 416412 7092
rect 416464 7080 416470 7132
rect 126974 7012 126980 7064
rect 127032 7052 127038 7064
rect 284294 7052 284300 7064
rect 127032 7024 284300 7052
rect 127032 7012 127038 7024
rect 284294 7012 284300 7024
rect 284352 7012 284358 7064
rect 355962 7012 355968 7064
rect 356020 7052 356026 7064
rect 403618 7052 403624 7064
rect 356020 7024 403624 7052
rect 356020 7012 356026 7024
rect 403618 7012 403624 7024
rect 403676 7012 403682 7064
rect 279510 6808 279516 6860
rect 279568 6848 279574 6860
rect 322934 6848 322940 6860
rect 279568 6820 322940 6848
rect 279568 6808 279574 6820
rect 322934 6808 322940 6820
rect 322992 6808 322998 6860
rect 350442 6808 350448 6860
rect 350500 6848 350506 6860
rect 382366 6848 382372 6860
rect 350500 6820 382372 6848
rect 350500 6808 350506 6820
rect 382366 6808 382372 6820
rect 382424 6808 382430 6860
rect 522298 6808 522304 6860
rect 522356 6848 522362 6860
rect 580166 6848 580172 6860
rect 522356 6820 580172 6848
rect 522356 6808 522362 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 209682 6740 209688 6792
rect 209740 6780 209746 6792
rect 285398 6780 285404 6792
rect 209740 6752 285404 6780
rect 209740 6740 209746 6752
rect 285398 6740 285404 6752
rect 285456 6740 285462 6792
rect 286594 6740 286600 6792
rect 286652 6780 286658 6792
rect 324314 6780 324320 6792
rect 286652 6752 324320 6780
rect 286652 6740 286658 6752
rect 324314 6740 324320 6752
rect 324372 6740 324378 6792
rect 325602 6740 325608 6792
rect 325660 6780 325666 6792
rect 335446 6780 335452 6792
rect 325660 6752 335452 6780
rect 325660 6740 325666 6752
rect 335446 6740 335452 6752
rect 335504 6740 335510 6792
rect 351730 6740 351736 6792
rect 351788 6780 351794 6792
rect 385954 6780 385960 6792
rect 351788 6752 385960 6780
rect 351788 6740 351794 6752
rect 385954 6740 385960 6752
rect 386012 6740 386018 6792
rect 391842 6740 391848 6792
rect 391900 6780 391906 6792
rect 545482 6780 545488 6792
rect 391900 6752 545488 6780
rect 391900 6740 391906 6752
rect 545482 6740 545488 6752
rect 545540 6740 545546 6792
rect 220078 6672 220084 6724
rect 220136 6712 220142 6724
rect 296070 6712 296076 6724
rect 220136 6684 296076 6712
rect 220136 6672 220142 6684
rect 296070 6672 296076 6684
rect 296128 6672 296134 6724
rect 297266 6672 297272 6724
rect 297324 6712 297330 6724
rect 327258 6712 327264 6724
rect 297324 6684 327264 6712
rect 297324 6672 297330 6684
rect 327258 6672 327264 6684
rect 327316 6672 327322 6724
rect 351822 6672 351828 6724
rect 351880 6712 351886 6724
rect 389450 6712 389456 6724
rect 351880 6684 389456 6712
rect 351880 6672 351886 6684
rect 389450 6672 389456 6684
rect 389508 6672 389514 6724
rect 393222 6672 393228 6724
rect 393280 6712 393286 6724
rect 549070 6712 549076 6724
rect 393280 6684 549076 6712
rect 393280 6672 393286 6684
rect 549070 6672 549076 6684
rect 549128 6672 549134 6724
rect 190822 6604 190828 6656
rect 190880 6644 190886 6656
rect 287698 6644 287704 6656
rect 190880 6616 287704 6644
rect 190880 6604 190886 6616
rect 287698 6604 287704 6616
rect 287756 6604 287762 6656
rect 290182 6604 290188 6656
rect 290240 6644 290246 6656
rect 325694 6644 325700 6656
rect 290240 6616 325700 6644
rect 290240 6604 290246 6616
rect 325694 6604 325700 6616
rect 325752 6604 325758 6656
rect 342162 6604 342168 6656
rect 342220 6644 342226 6656
rect 350442 6644 350448 6656
rect 342220 6616 350448 6644
rect 342220 6604 342226 6616
rect 350442 6604 350448 6616
rect 350500 6604 350506 6656
rect 353202 6604 353208 6656
rect 353260 6644 353266 6656
rect 393038 6644 393044 6656
rect 353260 6616 393044 6644
rect 353260 6604 353266 6616
rect 393038 6604 393044 6616
rect 393096 6604 393102 6656
rect 394510 6604 394516 6656
rect 394568 6644 394574 6656
rect 552658 6644 552664 6656
rect 394568 6616 552664 6644
rect 394568 6604 394574 6616
rect 552658 6604 552664 6616
rect 552716 6604 552722 6656
rect 176654 6536 176660 6588
rect 176712 6576 176718 6588
rect 291838 6576 291844 6588
rect 176712 6548 291844 6576
rect 176712 6536 176718 6548
rect 291838 6536 291844 6548
rect 291896 6536 291902 6588
rect 293678 6536 293684 6588
rect 293736 6576 293742 6588
rect 327166 6576 327172 6588
rect 293736 6548 327172 6576
rect 293736 6536 293742 6548
rect 327166 6536 327172 6548
rect 327224 6536 327230 6588
rect 343542 6536 343548 6588
rect 343600 6576 343606 6588
rect 354030 6576 354036 6588
rect 343600 6548 354036 6576
rect 343600 6536 343606 6548
rect 354030 6536 354036 6548
rect 354088 6536 354094 6588
rect 354582 6536 354588 6588
rect 354640 6576 354646 6588
rect 354640 6548 393314 6576
rect 354640 6536 354646 6548
rect 230290 6468 230296 6520
rect 230348 6508 230354 6520
rect 363506 6508 363512 6520
rect 230348 6480 363512 6508
rect 230348 6468 230354 6480
rect 363506 6468 363512 6480
rect 363564 6468 363570 6520
rect 230382 6400 230388 6452
rect 230440 6440 230446 6452
rect 367002 6440 367008 6452
rect 230440 6412 367008 6440
rect 230440 6400 230446 6412
rect 367002 6400 367008 6412
rect 367060 6400 367066 6452
rect 393286 6440 393314 6548
rect 394602 6536 394608 6588
rect 394660 6576 394666 6588
rect 556154 6576 556160 6588
rect 394660 6548 556160 6576
rect 394660 6536 394666 6548
rect 556154 6536 556160 6548
rect 556212 6536 556218 6588
rect 395890 6468 395896 6520
rect 395948 6508 395954 6520
rect 559742 6508 559748 6520
rect 395948 6480 559748 6508
rect 395948 6468 395954 6480
rect 559742 6468 559748 6480
rect 559800 6468 559806 6520
rect 396534 6440 396540 6452
rect 393286 6412 396540 6440
rect 396534 6400 396540 6412
rect 396592 6400 396598 6452
rect 397362 6400 397368 6452
rect 397420 6440 397426 6452
rect 563238 6440 563244 6452
rect 397420 6412 563244 6440
rect 397420 6400 397426 6412
rect 563238 6400 563244 6412
rect 563296 6400 563302 6452
rect 231762 6332 231768 6384
rect 231820 6372 231826 6384
rect 370590 6372 370596 6384
rect 231820 6344 370596 6372
rect 231820 6332 231826 6344
rect 370590 6332 370596 6344
rect 370648 6332 370654 6384
rect 397270 6332 397276 6384
rect 397328 6372 397334 6384
rect 566826 6372 566832 6384
rect 397328 6344 566832 6372
rect 397328 6332 397334 6344
rect 566826 6332 566832 6344
rect 566884 6332 566890 6384
rect 233050 6264 233056 6316
rect 233108 6304 233114 6316
rect 374086 6304 374092 6316
rect 233108 6276 374092 6304
rect 233108 6264 233114 6276
rect 374086 6264 374092 6276
rect 374144 6264 374150 6316
rect 374638 6264 374644 6316
rect 374696 6304 374702 6316
rect 384758 6304 384764 6316
rect 374696 6276 384764 6304
rect 374696 6264 374702 6276
rect 384758 6264 384764 6276
rect 384816 6264 384822 6316
rect 398742 6264 398748 6316
rect 398800 6304 398806 6316
rect 570322 6304 570328 6316
rect 398800 6276 570328 6304
rect 398800 6264 398806 6276
rect 570322 6264 570328 6276
rect 570380 6264 570386 6316
rect 233142 6196 233148 6248
rect 233200 6236 233206 6248
rect 377674 6236 377680 6248
rect 233200 6208 377680 6236
rect 233200 6196 233206 6208
rect 377674 6196 377680 6208
rect 377732 6196 377738 6248
rect 391750 6196 391756 6248
rect 391808 6236 391814 6248
rect 398101 6239 398159 6245
rect 398101 6236 398113 6239
rect 391808 6208 398113 6236
rect 391808 6196 391814 6208
rect 398101 6205 398113 6208
rect 398147 6205 398159 6239
rect 398101 6199 398159 6205
rect 400122 6196 400128 6248
rect 400180 6236 400186 6248
rect 573910 6236 573916 6248
rect 400180 6208 573916 6236
rect 400180 6196 400186 6208
rect 573910 6196 573916 6208
rect 573968 6196 573974 6248
rect 234522 6128 234528 6180
rect 234580 6168 234586 6180
rect 381170 6168 381176 6180
rect 234580 6140 381176 6168
rect 234580 6128 234586 6140
rect 381170 6128 381176 6140
rect 381228 6128 381234 6180
rect 384850 6128 384856 6180
rect 384908 6168 384914 6180
rect 391937 6171 391995 6177
rect 391937 6168 391949 6171
rect 384908 6140 391949 6168
rect 384908 6128 384914 6140
rect 391937 6137 391949 6140
rect 391983 6137 391995 6171
rect 391937 6131 391995 6137
rect 398009 6171 398067 6177
rect 398009 6137 398021 6171
rect 398055 6168 398067 6171
rect 399938 6168 399944 6180
rect 398055 6140 399944 6168
rect 398055 6137 398067 6140
rect 398009 6131 398067 6137
rect 399938 6128 399944 6140
rect 399996 6128 400002 6180
rect 400030 6128 400036 6180
rect 400088 6168 400094 6180
rect 577406 6168 577412 6180
rect 400088 6140 577412 6168
rect 400088 6128 400094 6140
rect 577406 6128 577412 6140
rect 577464 6128 577470 6180
rect 272426 6060 272432 6112
rect 272484 6100 272490 6112
rect 305638 6100 305644 6112
rect 272484 6072 305644 6100
rect 272484 6060 272490 6072
rect 305638 6060 305644 6072
rect 305696 6060 305702 6112
rect 307938 6060 307944 6112
rect 307996 6100 308002 6112
rect 329926 6100 329932 6112
rect 307996 6072 329932 6100
rect 307996 6060 308002 6072
rect 329926 6060 329932 6072
rect 329984 6060 329990 6112
rect 349062 6060 349068 6112
rect 349120 6100 349126 6112
rect 378870 6100 378876 6112
rect 349120 6072 378876 6100
rect 349120 6060 349126 6072
rect 378870 6060 378876 6072
rect 378928 6060 378934 6112
rect 390462 6060 390468 6112
rect 390520 6100 390526 6112
rect 538398 6100 538404 6112
rect 390520 6072 538404 6100
rect 390520 6060 390526 6072
rect 538398 6060 538404 6072
rect 538456 6060 538462 6112
rect 264238 5992 264244 6044
rect 264296 6032 264302 6044
rect 292574 6032 292580 6044
rect 264296 6004 292580 6032
rect 264296 5992 264302 6004
rect 292574 5992 292580 6004
rect 292632 5992 292638 6044
rect 300762 5992 300768 6044
rect 300820 6032 300826 6044
rect 328454 6032 328460 6044
rect 300820 6004 328460 6032
rect 300820 5992 300826 6004
rect 328454 5992 328460 6004
rect 328512 5992 328518 6044
rect 348970 5992 348976 6044
rect 349028 6032 349034 6044
rect 375282 6032 375288 6044
rect 349028 6004 375288 6032
rect 349028 5992 349034 6004
rect 375282 5992 375288 6004
rect 375340 5992 375346 6044
rect 389082 5992 389088 6044
rect 389140 6032 389146 6044
rect 534902 6032 534908 6044
rect 389140 6004 534908 6032
rect 389140 5992 389146 6004
rect 534902 5992 534908 6004
rect 534960 5992 534966 6044
rect 265342 5924 265348 5976
rect 265400 5964 265406 5976
rect 286318 5964 286324 5976
rect 265400 5936 286324 5964
rect 265400 5924 265406 5936
rect 286318 5924 286324 5936
rect 286376 5924 286382 5976
rect 304350 5924 304356 5976
rect 304408 5964 304414 5976
rect 329834 5964 329840 5976
rect 304408 5936 329840 5964
rect 304408 5924 304414 5936
rect 329834 5924 329840 5936
rect 329892 5924 329898 5976
rect 347682 5924 347688 5976
rect 347740 5964 347746 5976
rect 371694 5964 371700 5976
rect 347740 5936 371700 5964
rect 347740 5924 347746 5936
rect 371694 5924 371700 5936
rect 371752 5924 371758 5976
rect 388990 5924 388996 5976
rect 389048 5964 389054 5976
rect 531314 5964 531320 5976
rect 389048 5936 531320 5964
rect 389048 5924 389054 5936
rect 531314 5924 531320 5936
rect 531372 5924 531378 5976
rect 311434 5856 311440 5908
rect 311492 5896 311498 5908
rect 331306 5896 331312 5908
rect 311492 5868 331312 5896
rect 311492 5856 311498 5868
rect 331306 5856 331312 5868
rect 331364 5856 331370 5908
rect 344830 5856 344836 5908
rect 344888 5896 344894 5908
rect 349893 5899 349951 5905
rect 349893 5896 349905 5899
rect 344888 5868 349905 5896
rect 344888 5856 344894 5868
rect 349893 5865 349905 5868
rect 349939 5865 349951 5899
rect 368198 5896 368204 5908
rect 349893 5859 349951 5865
rect 350000 5868 368204 5896
rect 315022 5788 315028 5840
rect 315080 5828 315086 5840
rect 332686 5828 332692 5840
rect 315080 5800 332692 5828
rect 315080 5788 315086 5800
rect 332686 5788 332692 5800
rect 332744 5788 332750 5840
rect 347590 5788 347596 5840
rect 347648 5828 347654 5840
rect 350000 5828 350028 5868
rect 368198 5856 368204 5868
rect 368256 5856 368262 5908
rect 387702 5856 387708 5908
rect 387760 5896 387766 5908
rect 527818 5896 527824 5908
rect 387760 5868 527824 5896
rect 387760 5856 387766 5868
rect 527818 5856 527824 5868
rect 527876 5856 527882 5908
rect 347648 5800 350028 5828
rect 350077 5831 350135 5837
rect 347648 5788 347654 5800
rect 350077 5797 350089 5831
rect 350123 5828 350135 5831
rect 364610 5828 364616 5840
rect 350123 5800 364616 5828
rect 350123 5797 350135 5800
rect 350077 5791 350135 5797
rect 364610 5788 364616 5800
rect 364668 5788 364674 5840
rect 386230 5788 386236 5840
rect 386288 5828 386294 5840
rect 524230 5828 524236 5840
rect 386288 5800 524236 5828
rect 386288 5788 386294 5800
rect 524230 5788 524236 5800
rect 524288 5788 524294 5840
rect 318518 5720 318524 5772
rect 318576 5760 318582 5772
rect 332594 5760 332600 5772
rect 318576 5732 332600 5760
rect 318576 5720 318582 5732
rect 332594 5720 332600 5732
rect 332652 5720 332658 5772
rect 344922 5720 344928 5772
rect 344980 5760 344986 5772
rect 349893 5763 349951 5769
rect 344980 5732 349844 5760
rect 344980 5720 344986 5732
rect 322106 5652 322112 5704
rect 322164 5692 322170 5704
rect 333974 5692 333980 5704
rect 322164 5664 333980 5692
rect 322164 5652 322170 5664
rect 333974 5652 333980 5664
rect 334032 5652 334038 5704
rect 342070 5652 342076 5704
rect 342128 5692 342134 5704
rect 346946 5692 346952 5704
rect 342128 5664 346952 5692
rect 342128 5652 342134 5664
rect 346946 5652 346952 5664
rect 347004 5652 347010 5704
rect 349816 5692 349844 5732
rect 349893 5729 349905 5763
rect 349939 5760 349951 5763
rect 361114 5760 361120 5772
rect 349939 5732 361120 5760
rect 349939 5729 349951 5732
rect 349893 5723 349951 5729
rect 361114 5720 361120 5732
rect 361172 5720 361178 5772
rect 386322 5720 386328 5772
rect 386380 5760 386386 5772
rect 520734 5760 520740 5772
rect 386380 5732 520740 5760
rect 386380 5720 386386 5732
rect 520734 5720 520740 5732
rect 520792 5720 520798 5772
rect 357526 5692 357532 5704
rect 349816 5664 357532 5692
rect 357526 5652 357532 5664
rect 357584 5652 357590 5704
rect 384942 5652 384948 5704
rect 385000 5692 385006 5704
rect 517146 5692 517152 5704
rect 385000 5664 517152 5692
rect 385000 5652 385006 5664
rect 517146 5652 517152 5664
rect 517204 5652 517210 5704
rect 329190 5584 329196 5636
rect 329248 5624 329254 5636
rect 335354 5624 335360 5636
rect 329248 5596 335360 5624
rect 329248 5584 329254 5596
rect 335354 5584 335360 5596
rect 335412 5584 335418 5636
rect 336734 5624 336740 5636
rect 336016 5596 336740 5624
rect 332686 5516 332692 5568
rect 332744 5556 332750 5568
rect 336016 5556 336044 5596
rect 336734 5584 336740 5596
rect 336792 5584 336798 5636
rect 346302 5584 346308 5636
rect 346360 5624 346366 5636
rect 350077 5627 350135 5633
rect 350077 5624 350089 5627
rect 346360 5596 350089 5624
rect 346360 5584 346366 5596
rect 350077 5593 350089 5596
rect 350123 5593 350135 5627
rect 350077 5587 350135 5593
rect 389818 5584 389824 5636
rect 389876 5624 389882 5636
rect 391842 5624 391848 5636
rect 389876 5596 391848 5624
rect 389876 5584 389882 5596
rect 391842 5584 391848 5596
rect 391900 5584 391906 5636
rect 391937 5627 391995 5633
rect 391937 5593 391949 5627
rect 391983 5624 391995 5627
rect 513558 5624 513564 5636
rect 391983 5596 513564 5624
rect 391983 5593 391995 5596
rect 391937 5587 391995 5593
rect 513558 5584 513564 5596
rect 513616 5584 513622 5636
rect 332744 5528 336044 5556
rect 332744 5516 332750 5528
rect 336274 5516 336280 5568
rect 336332 5556 336338 5568
rect 338114 5556 338120 5568
rect 336332 5528 338120 5556
rect 336332 5516 336338 5528
rect 338114 5516 338120 5528
rect 338172 5516 338178 5568
rect 339402 5516 339408 5568
rect 339460 5556 339466 5568
rect 339862 5556 339868 5568
rect 339460 5528 339868 5556
rect 339460 5516 339466 5528
rect 339862 5516 339868 5528
rect 339920 5516 339926 5568
rect 340782 5516 340788 5568
rect 340840 5556 340846 5568
rect 343358 5556 343364 5568
rect 340840 5528 343364 5556
rect 340840 5516 340846 5528
rect 343358 5516 343364 5528
rect 343416 5516 343422 5568
rect 354490 5516 354496 5568
rect 354548 5556 354554 5568
rect 398009 5559 398067 5565
rect 398009 5556 398021 5559
rect 354548 5528 398021 5556
rect 354548 5516 354554 5528
rect 398009 5525 398021 5528
rect 398055 5525 398067 5559
rect 398009 5519 398067 5525
rect 398101 5559 398159 5565
rect 398101 5525 398113 5559
rect 398147 5556 398159 5559
rect 541986 5556 541992 5568
rect 398147 5528 541992 5556
rect 398147 5525 398159 5528
rect 398101 5519 398159 5525
rect 541986 5516 541992 5528
rect 542044 5516 542050 5568
rect 200022 5448 200028 5500
rect 200080 5488 200086 5500
rect 246390 5488 246396 5500
rect 200080 5460 246396 5488
rect 200080 5448 200086 5460
rect 246390 5448 246396 5460
rect 246448 5448 246454 5500
rect 274450 5448 274456 5500
rect 274508 5488 274514 5500
rect 540790 5488 540796 5500
rect 274508 5460 540796 5488
rect 274508 5448 274514 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 201310 5380 201316 5432
rect 201368 5420 201374 5432
rect 249978 5420 249984 5432
rect 201368 5392 249984 5420
rect 201368 5380 201374 5392
rect 249978 5380 249984 5392
rect 250036 5380 250042 5432
rect 275922 5380 275928 5432
rect 275980 5420 275986 5432
rect 544378 5420 544384 5432
rect 275980 5392 544384 5420
rect 275980 5380 275986 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 201402 5312 201408 5364
rect 201460 5352 201466 5364
rect 253474 5352 253480 5364
rect 201460 5324 253480 5352
rect 201460 5312 201466 5324
rect 253474 5312 253480 5324
rect 253532 5312 253538 5364
rect 277302 5312 277308 5364
rect 277360 5352 277366 5364
rect 547874 5352 547880 5364
rect 277360 5324 547880 5352
rect 277360 5312 277366 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 202782 5244 202788 5296
rect 202840 5284 202846 5296
rect 257062 5284 257068 5296
rect 202840 5256 257068 5284
rect 202840 5244 202846 5256
rect 257062 5244 257068 5256
rect 257120 5244 257126 5296
rect 277210 5244 277216 5296
rect 277268 5284 277274 5296
rect 551462 5284 551468 5296
rect 277268 5256 551468 5284
rect 277268 5244 277274 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 202690 5176 202696 5228
rect 202748 5216 202754 5228
rect 260558 5216 260564 5228
rect 202748 5188 260564 5216
rect 202748 5176 202754 5188
rect 260558 5176 260564 5188
rect 260616 5176 260622 5228
rect 278682 5176 278688 5228
rect 278740 5216 278746 5228
rect 554958 5216 554964 5228
rect 278740 5188 554964 5216
rect 278740 5176 278746 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 204162 5108 204168 5160
rect 204220 5148 204226 5160
rect 264146 5148 264152 5160
rect 204220 5120 264152 5148
rect 204220 5108 204226 5120
rect 264146 5108 264152 5120
rect 264204 5108 264210 5160
rect 279970 5108 279976 5160
rect 280028 5148 280034 5160
rect 558546 5148 558552 5160
rect 280028 5120 558552 5148
rect 280028 5108 280034 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 205542 5040 205548 5092
rect 205600 5080 205606 5092
rect 267734 5080 267740 5092
rect 205600 5052 267740 5080
rect 205600 5040 205606 5052
rect 267734 5040 267740 5052
rect 267792 5040 267798 5092
rect 280062 5040 280068 5092
rect 280120 5080 280126 5092
rect 562042 5080 562048 5092
rect 280120 5052 562048 5080
rect 280120 5040 280126 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 205450 4972 205456 5024
rect 205508 5012 205514 5024
rect 271230 5012 271236 5024
rect 205508 4984 271236 5012
rect 205508 4972 205514 4984
rect 271230 4972 271236 4984
rect 271288 4972 271294 5024
rect 281442 4972 281448 5024
rect 281500 5012 281506 5024
rect 565630 5012 565636 5024
rect 281500 4984 565636 5012
rect 281500 4972 281506 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 206922 4904 206928 4956
rect 206980 4944 206986 4956
rect 274818 4944 274824 4956
rect 206980 4916 274824 4944
rect 206980 4904 206986 4916
rect 274818 4904 274824 4916
rect 274876 4904 274882 4956
rect 282822 4904 282828 4956
rect 282880 4944 282886 4956
rect 569126 4944 569132 4956
rect 282880 4916 569132 4944
rect 282880 4904 282886 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 208210 4836 208216 4888
rect 208268 4876 208274 4888
rect 278314 4876 278320 4888
rect 208268 4848 278320 4876
rect 208268 4836 208274 4848
rect 278314 4836 278320 4848
rect 278372 4836 278378 4888
rect 282730 4836 282736 4888
rect 282788 4876 282794 4888
rect 572714 4876 572720 4888
rect 282788 4848 572720 4876
rect 282788 4836 282794 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 208302 4768 208308 4820
rect 208360 4808 208366 4820
rect 281902 4808 281908 4820
rect 208360 4780 281908 4808
rect 208360 4768 208366 4780
rect 281902 4768 281908 4780
rect 281960 4768 281966 4820
rect 284202 4768 284208 4820
rect 284260 4808 284266 4820
rect 576302 4808 576308 4820
rect 284260 4780 576308 4808
rect 284260 4768 284266 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 198550 4700 198556 4752
rect 198608 4740 198614 4752
rect 242894 4740 242900 4752
rect 198608 4712 242900 4740
rect 198608 4700 198614 4712
rect 242894 4700 242900 4712
rect 242952 4700 242958 4752
rect 274542 4700 274548 4752
rect 274600 4740 274606 4752
rect 537202 4740 537208 4752
rect 274600 4712 537208 4740
rect 274600 4700 274606 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 198642 4632 198648 4684
rect 198700 4672 198706 4684
rect 239306 4672 239312 4684
rect 198700 4644 239312 4672
rect 198700 4632 198706 4644
rect 239306 4632 239312 4644
rect 239364 4632 239370 4684
rect 273070 4632 273076 4684
rect 273128 4672 273134 4684
rect 533706 4672 533712 4684
rect 273128 4644 533712 4672
rect 273128 4632 273134 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 197262 4564 197268 4616
rect 197320 4604 197326 4616
rect 235810 4604 235816 4616
rect 197320 4576 235816 4604
rect 197320 4564 197326 4576
rect 235810 4564 235816 4576
rect 235868 4564 235874 4616
rect 273162 4564 273168 4616
rect 273220 4604 273226 4616
rect 530118 4604 530124 4616
rect 273220 4576 530124 4604
rect 273220 4564 273226 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 195790 4496 195796 4548
rect 195848 4536 195854 4548
rect 232222 4536 232228 4548
rect 195848 4508 232228 4536
rect 195848 4496 195854 4508
rect 232222 4496 232228 4508
rect 232280 4496 232286 4548
rect 271782 4496 271788 4548
rect 271840 4536 271846 4548
rect 526622 4536 526628 4548
rect 271840 4508 526628 4536
rect 271840 4496 271846 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 195882 4428 195888 4480
rect 195940 4468 195946 4480
rect 228726 4468 228732 4480
rect 195940 4440 228732 4468
rect 195940 4428 195946 4440
rect 228726 4428 228732 4440
rect 228784 4428 228790 4480
rect 270402 4428 270408 4480
rect 270460 4468 270466 4480
rect 523034 4468 523040 4480
rect 270460 4440 523040 4468
rect 270460 4428 270466 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 194502 4360 194508 4412
rect 194560 4400 194566 4412
rect 225138 4400 225144 4412
rect 194560 4372 225144 4400
rect 194560 4360 194566 4372
rect 225138 4360 225144 4372
rect 225196 4360 225202 4412
rect 270310 4360 270316 4412
rect 270368 4400 270374 4412
rect 519538 4400 519544 4412
rect 270368 4372 519544 4400
rect 270368 4360 270374 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 193122 4292 193128 4344
rect 193180 4332 193186 4344
rect 221550 4332 221556 4344
rect 193180 4304 221556 4332
rect 193180 4292 193186 4304
rect 221550 4292 221556 4304
rect 221608 4292 221614 4344
rect 269022 4292 269028 4344
rect 269080 4332 269086 4344
rect 515950 4332 515956 4344
rect 269080 4304 515956 4332
rect 269080 4292 269086 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 193030 4224 193036 4276
rect 193088 4264 193094 4276
rect 218054 4264 218060 4276
rect 193088 4236 218060 4264
rect 193088 4224 193094 4236
rect 218054 4224 218060 4236
rect 218112 4224 218118 4276
rect 267642 4224 267648 4276
rect 267700 4264 267706 4276
rect 512454 4264 512460 4276
rect 267700 4236 512460 4264
rect 267700 4224 267706 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 400858 4156 400864 4208
rect 400916 4196 400922 4208
rect 402514 4196 402520 4208
rect 400916 4168 402520 4196
rect 400916 4156 400922 4168
rect 402514 4156 402520 4168
rect 402572 4156 402578 4208
rect 454405 4199 454463 4205
rect 454405 4165 454417 4199
rect 454451 4196 454463 4199
rect 456794 4196 456800 4208
rect 454451 4168 456800 4196
rect 454451 4165 454463 4168
rect 454405 4159 454463 4165
rect 456794 4156 456800 4168
rect 456852 4156 456858 4208
rect 340966 4088 340972 4140
rect 341024 4128 341030 4140
rect 377398 4128 377404 4140
rect 341024 4100 377404 4128
rect 341024 4088 341030 4100
rect 377398 4088 377404 4100
rect 377456 4088 377462 4140
rect 394234 4088 394240 4140
rect 394292 4128 394298 4140
rect 467834 4128 467840 4140
rect 394292 4100 467840 4128
rect 394292 4088 394298 4100
rect 467834 4088 467840 4100
rect 467892 4088 467898 4140
rect 507762 4088 507768 4140
rect 507820 4128 507826 4140
rect 543182 4128 543188 4140
rect 507820 4100 543188 4128
rect 507820 4088 507826 4100
rect 543182 4088 543188 4100
rect 543240 4088 543246 4140
rect 319714 4020 319720 4072
rect 319772 4060 319778 4072
rect 356698 4060 356704 4072
rect 319772 4032 356704 4060
rect 319772 4020 319778 4032
rect 356698 4020 356704 4032
rect 356756 4020 356762 4072
rect 390646 4020 390652 4072
rect 390704 4060 390710 4072
rect 461029 4063 461087 4069
rect 461029 4060 461041 4063
rect 390704 4032 461041 4060
rect 390704 4020 390710 4032
rect 461029 4029 461041 4032
rect 461075 4029 461087 4063
rect 466454 4060 466460 4072
rect 461029 4023 461087 4029
rect 461136 4032 466460 4060
rect 138842 3952 138848 4004
rect 138900 3992 138906 4004
rect 142798 3992 142804 4004
rect 138900 3964 142804 3992
rect 138900 3952 138906 3964
rect 142798 3952 142804 3964
rect 142856 3952 142862 4004
rect 196618 3952 196624 4004
rect 196676 3992 196682 4004
rect 203886 3992 203892 4004
rect 196676 3964 203892 3992
rect 196676 3952 196682 3964
rect 203886 3952 203892 3964
rect 203944 3952 203950 4004
rect 309042 3952 309048 4004
rect 309100 3992 309106 4004
rect 340138 3992 340144 4004
rect 309100 3964 340144 3992
rect 309100 3952 309106 3964
rect 340138 3952 340144 3964
rect 340196 3952 340202 4004
rect 344554 3952 344560 4004
rect 344612 3992 344618 4004
rect 382918 3992 382924 4004
rect 344612 3964 382924 3992
rect 344612 3952 344618 3964
rect 382918 3952 382924 3964
rect 382976 3952 382982 4004
rect 387150 3952 387156 4004
rect 387208 3992 387214 4004
rect 461136 3992 461164 4032
rect 466454 4020 466460 4032
rect 466512 4020 466518 4072
rect 489178 4020 489184 4072
rect 489236 4060 489242 4072
rect 491110 4060 491116 4072
rect 489236 4032 491116 4060
rect 489236 4020 489242 4032
rect 491110 4020 491116 4032
rect 491168 4020 491174 4072
rect 509050 4020 509056 4072
rect 509108 4060 509114 4072
rect 546678 4060 546684 4072
rect 509108 4032 546684 4060
rect 509108 4020 509114 4032
rect 546678 4020 546684 4032
rect 546736 4020 546742 4072
rect 387208 3964 461164 3992
rect 461213 3995 461271 4001
rect 387208 3952 387214 3964
rect 461213 3961 461225 3995
rect 461259 3992 461271 3995
rect 465166 3992 465172 4004
rect 461259 3964 465172 3992
rect 461259 3961 461271 3964
rect 461213 3955 461271 3961
rect 465166 3952 465172 3964
rect 465224 3952 465230 4004
rect 497458 3952 497464 4004
rect 497516 3992 497522 4004
rect 500586 3992 500592 4004
rect 497516 3964 500592 3992
rect 497516 3952 497522 3964
rect 500586 3952 500592 3964
rect 500644 3952 500650 4004
rect 509142 3952 509148 4004
rect 509200 3992 509206 4004
rect 550266 3992 550272 4004
rect 509200 3964 550272 3992
rect 509200 3952 509206 3964
rect 550266 3952 550272 3964
rect 550324 3952 550330 4004
rect 164789 3927 164847 3933
rect 164789 3893 164801 3927
rect 164835 3924 164847 3927
rect 169018 3924 169024 3936
rect 164835 3896 169024 3924
rect 164835 3893 164847 3896
rect 164789 3887 164847 3893
rect 169018 3884 169024 3896
rect 169076 3884 169082 3936
rect 187602 3884 187608 3936
rect 187660 3924 187666 3936
rect 196802 3924 196808 3936
rect 187660 3896 196808 3924
rect 187660 3884 187666 3896
rect 196802 3884 196808 3896
rect 196860 3884 196866 3936
rect 248782 3884 248788 3936
rect 248840 3924 248846 3936
rect 266998 3924 267004 3936
rect 248840 3896 267004 3924
rect 248840 3884 248846 3896
rect 266998 3884 267004 3896
rect 267056 3884 267062 3936
rect 277210 3884 277216 3936
rect 277268 3924 277274 3936
rect 294598 3924 294604 3936
rect 277268 3896 294604 3924
rect 277268 3884 277274 3896
rect 294598 3884 294604 3896
rect 294656 3884 294662 3936
rect 301958 3884 301964 3936
rect 302016 3924 302022 3936
rect 318058 3924 318064 3936
rect 302016 3896 318064 3924
rect 302016 3884 302022 3896
rect 318058 3884 318064 3896
rect 318116 3884 318122 3936
rect 326798 3884 326804 3936
rect 326856 3924 326862 3936
rect 363598 3924 363604 3936
rect 326856 3896 363604 3924
rect 326856 3884 326862 3896
rect 363598 3884 363604 3896
rect 363656 3884 363662 3936
rect 383562 3884 383568 3936
rect 383620 3924 383626 3936
rect 465258 3924 465264 3936
rect 383620 3896 465264 3924
rect 383620 3884 383626 3896
rect 465258 3884 465264 3896
rect 465316 3884 465322 3936
rect 511902 3884 511908 3936
rect 511960 3924 511966 3936
rect 515677 3927 515735 3933
rect 515677 3924 515689 3927
rect 511960 3896 515689 3924
rect 511960 3884 511966 3896
rect 515677 3893 515689 3896
rect 515723 3893 515735 3927
rect 515677 3887 515735 3893
rect 515769 3927 515827 3933
rect 515769 3893 515781 3927
rect 515815 3924 515827 3927
rect 553762 3924 553768 3936
rect 515815 3896 553768 3924
rect 515815 3893 515827 3896
rect 515769 3887 515827 3893
rect 553762 3884 553768 3896
rect 553820 3884 553826 3936
rect 154206 3816 154212 3868
rect 154264 3856 154270 3868
rect 166258 3856 166264 3868
rect 154264 3828 166264 3856
rect 154264 3816 154270 3828
rect 166258 3816 166264 3828
rect 166316 3816 166322 3868
rect 168374 3816 168380 3868
rect 168432 3856 168438 3868
rect 178218 3856 178224 3868
rect 168432 3828 178224 3856
rect 168432 3816 168438 3828
rect 178218 3816 178224 3828
rect 178276 3816 178282 3868
rect 190270 3816 190276 3868
rect 190328 3856 190334 3868
rect 207382 3856 207388 3868
rect 190328 3828 207388 3856
rect 190328 3816 190334 3828
rect 207382 3816 207388 3828
rect 207440 3816 207446 3868
rect 271138 3856 271144 3868
rect 258046 3828 271144 3856
rect 145926 3748 145932 3800
rect 145984 3788 145990 3800
rect 162118 3788 162124 3800
rect 145984 3760 162124 3788
rect 145984 3748 145990 3760
rect 162118 3748 162124 3760
rect 162176 3748 162182 3800
rect 166074 3748 166080 3800
rect 166132 3788 166138 3800
rect 177298 3788 177304 3800
rect 166132 3760 177304 3788
rect 166132 3748 166138 3760
rect 177298 3748 177304 3760
rect 177356 3748 177362 3800
rect 190362 3748 190368 3800
rect 190420 3788 190426 3800
rect 210970 3788 210976 3800
rect 190420 3760 210976 3788
rect 190420 3748 190426 3760
rect 210970 3748 210976 3760
rect 211028 3748 211034 3800
rect 252370 3748 252376 3800
rect 252428 3788 252434 3800
rect 258046 3788 258074 3828
rect 271138 3816 271144 3828
rect 271196 3816 271202 3868
rect 294874 3816 294880 3868
rect 294932 3856 294938 3868
rect 323578 3856 323584 3868
rect 294932 3828 323584 3856
rect 294932 3816 294938 3828
rect 323578 3816 323584 3828
rect 323636 3816 323642 3868
rect 337470 3816 337476 3868
rect 337528 3856 337534 3868
rect 376018 3856 376024 3868
rect 337528 3828 376024 3856
rect 337528 3816 337534 3828
rect 376018 3816 376024 3828
rect 376076 3816 376082 3868
rect 379974 3816 379980 3868
rect 380032 3856 380038 3868
rect 461213 3859 461271 3865
rect 461213 3856 461225 3859
rect 380032 3828 461225 3856
rect 380032 3816 380038 3828
rect 461213 3825 461225 3828
rect 461259 3825 461271 3859
rect 463694 3856 463700 3868
rect 461213 3819 461271 3825
rect 461320 3828 463700 3856
rect 252428 3760 258074 3788
rect 252428 3748 252434 3760
rect 266538 3748 266544 3800
rect 266596 3788 266602 3800
rect 295978 3788 295984 3800
rect 266596 3760 295984 3788
rect 266596 3748 266602 3760
rect 295978 3748 295984 3760
rect 296036 3748 296042 3800
rect 298462 3748 298468 3800
rect 298520 3788 298526 3800
rect 320818 3788 320824 3800
rect 298520 3760 320824 3788
rect 298520 3748 298526 3760
rect 320818 3748 320824 3760
rect 320876 3748 320882 3800
rect 323302 3748 323308 3800
rect 323360 3788 323366 3800
rect 360838 3788 360844 3800
rect 323360 3760 360844 3788
rect 323360 3748 323366 3760
rect 360838 3748 360844 3760
rect 360896 3748 360902 3800
rect 376478 3748 376484 3800
rect 376536 3788 376542 3800
rect 461320 3788 461348 3828
rect 463694 3816 463700 3828
rect 463752 3816 463758 3868
rect 511810 3816 511816 3868
rect 511868 3856 511874 3868
rect 557350 3856 557356 3868
rect 511868 3828 557356 3856
rect 511868 3816 511874 3828
rect 557350 3816 557356 3828
rect 557408 3816 557414 3868
rect 462406 3788 462412 3800
rect 376536 3760 461348 3788
rect 461412 3760 462412 3788
rect 376536 3748 376542 3760
rect 160094 3680 160100 3732
rect 160152 3720 160158 3732
rect 188338 3720 188344 3732
rect 160152 3692 188344 3720
rect 160152 3680 160158 3692
rect 188338 3680 188344 3692
rect 188396 3680 188402 3732
rect 191742 3680 191748 3732
rect 191800 3720 191806 3732
rect 214466 3720 214472 3732
rect 191800 3692 214472 3720
rect 191800 3680 191806 3692
rect 214466 3680 214472 3692
rect 214524 3680 214530 3732
rect 238110 3680 238116 3732
rect 238168 3720 238174 3732
rect 249058 3720 249064 3732
rect 238168 3692 249064 3720
rect 238168 3680 238174 3692
rect 249058 3680 249064 3692
rect 249116 3680 249122 3732
rect 255866 3680 255872 3732
rect 255924 3720 255930 3732
rect 280798 3720 280804 3732
rect 255924 3692 280804 3720
rect 255924 3680 255930 3692
rect 280798 3680 280804 3692
rect 280856 3680 280862 3732
rect 287790 3680 287796 3732
rect 287848 3720 287854 3732
rect 322198 3720 322204 3732
rect 287848 3692 322204 3720
rect 287848 3680 287854 3692
rect 322198 3680 322204 3692
rect 322256 3680 322262 3732
rect 330386 3680 330392 3732
rect 330444 3720 330450 3732
rect 371878 3720 371884 3732
rect 330444 3692 371884 3720
rect 330444 3680 330450 3692
rect 371878 3680 371884 3692
rect 371936 3680 371942 3732
rect 372890 3680 372896 3732
rect 372948 3720 372954 3732
rect 452473 3723 452531 3729
rect 452473 3720 452485 3723
rect 372948 3692 452485 3720
rect 372948 3680 372954 3692
rect 452473 3689 452485 3692
rect 452519 3689 452531 3723
rect 461412 3720 461440 3760
rect 462406 3748 462412 3760
rect 462464 3748 462470 3800
rect 462590 3748 462596 3800
rect 462648 3788 462654 3800
rect 469214 3788 469220 3800
rect 462648 3760 469220 3788
rect 462648 3748 462654 3760
rect 469214 3748 469220 3760
rect 469272 3748 469278 3800
rect 498102 3748 498108 3800
rect 498160 3788 498166 3800
rect 504174 3788 504180 3800
rect 498160 3760 504180 3788
rect 498160 3748 498166 3760
rect 504174 3748 504180 3760
rect 504232 3748 504238 3800
rect 513282 3748 513288 3800
rect 513340 3788 513346 3800
rect 515677 3791 515735 3797
rect 513340 3760 515628 3788
rect 513340 3748 513346 3760
rect 452473 3683 452531 3689
rect 452672 3692 461440 3720
rect 461489 3723 461547 3729
rect 153010 3612 153016 3664
rect 153068 3652 153074 3664
rect 173066 3652 173072 3664
rect 153068 3624 173072 3652
rect 153068 3612 153074 3624
rect 173066 3612 173072 3624
rect 173124 3612 173130 3664
rect 180242 3612 180248 3664
rect 180300 3652 180306 3664
rect 184198 3652 184204 3664
rect 180300 3624 184204 3652
rect 180300 3612 180306 3624
rect 184198 3612 184204 3624
rect 184256 3612 184262 3664
rect 184308 3624 186268 3652
rect 137646 3544 137652 3596
rect 137704 3584 137710 3596
rect 164789 3587 164847 3593
rect 164789 3584 164801 3587
rect 137704 3556 164801 3584
rect 137704 3544 137710 3556
rect 164789 3553 164801 3556
rect 164835 3553 164847 3587
rect 164789 3547 164847 3553
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 165522 3584 165528 3596
rect 164936 3556 165528 3584
rect 164936 3544 164942 3556
rect 165522 3544 165528 3556
rect 165580 3544 165586 3596
rect 167178 3544 167184 3596
rect 167236 3584 167242 3596
rect 168282 3584 168288 3596
rect 167236 3556 168288 3584
rect 167236 3544 167242 3556
rect 168282 3544 168288 3556
rect 168340 3544 168346 3596
rect 173158 3544 173164 3596
rect 173216 3584 173222 3596
rect 173802 3584 173808 3596
rect 173216 3556 173808 3584
rect 173216 3544 173222 3556
rect 173802 3544 173808 3556
rect 173860 3544 173866 3596
rect 179046 3544 179052 3596
rect 179104 3584 179110 3596
rect 180058 3584 180064 3596
rect 179104 3556 180064 3584
rect 179104 3544 179110 3556
rect 180058 3544 180064 3556
rect 180116 3544 180122 3596
rect 181438 3544 181444 3596
rect 181496 3584 181502 3596
rect 182082 3584 182088 3596
rect 181496 3556 182088 3584
rect 181496 3544 181502 3556
rect 182082 3544 182088 3556
rect 182140 3544 182146 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 184308 3584 184336 3624
rect 183796 3556 184336 3584
rect 183796 3544 183802 3556
rect 184842 3544 184848 3596
rect 184900 3584 184906 3596
rect 186130 3584 186136 3596
rect 184900 3556 186136 3584
rect 184900 3544 184906 3556
rect 186130 3544 186136 3556
rect 186188 3544 186194 3596
rect 186240 3584 186268 3624
rect 187326 3612 187332 3664
rect 187384 3652 187390 3664
rect 214558 3652 214564 3664
rect 187384 3624 214564 3652
rect 187384 3612 187390 3624
rect 214558 3612 214564 3624
rect 214616 3612 214622 3664
rect 220446 3612 220452 3664
rect 220504 3652 220510 3664
rect 238018 3652 238024 3664
rect 220504 3624 238024 3652
rect 220504 3612 220510 3624
rect 238018 3612 238024 3624
rect 238076 3612 238082 3664
rect 260098 3652 260104 3664
rect 258046 3624 260104 3652
rect 224218 3584 224224 3596
rect 186240 3556 224224 3584
rect 224218 3544 224224 3556
rect 224276 3544 224282 3596
rect 231026 3544 231032 3596
rect 231084 3584 231090 3596
rect 231670 3584 231676 3596
rect 231084 3556 231676 3584
rect 231084 3544 231090 3556
rect 231670 3544 231676 3556
rect 231728 3544 231734 3596
rect 234614 3544 234620 3596
rect 234672 3584 234678 3596
rect 258046 3584 258074 3624
rect 260098 3612 260104 3624
rect 260156 3612 260162 3664
rect 262950 3612 262956 3664
rect 263008 3652 263014 3664
rect 298830 3652 298836 3664
rect 263008 3624 298836 3652
rect 263008 3612 263014 3624
rect 298830 3612 298836 3624
rect 298888 3612 298894 3664
rect 316218 3612 316224 3664
rect 316276 3652 316282 3664
rect 358078 3652 358084 3664
rect 316276 3624 358084 3652
rect 316276 3612 316282 3624
rect 358078 3612 358084 3624
rect 358136 3612 358142 3664
rect 369394 3612 369400 3664
rect 369452 3652 369458 3664
rect 452672 3652 452700 3692
rect 461489 3689 461501 3723
rect 461535 3720 461547 3723
rect 472066 3720 472072 3732
rect 461535 3692 472072 3720
rect 461535 3689 461547 3692
rect 461489 3683 461547 3689
rect 472066 3680 472072 3692
rect 472124 3680 472130 3732
rect 483750 3680 483756 3732
rect 483808 3720 483814 3732
rect 487157 3723 487215 3729
rect 487157 3720 487169 3723
rect 483808 3692 487169 3720
rect 483808 3680 483814 3692
rect 487157 3689 487169 3692
rect 487203 3689 487215 3723
rect 487157 3683 487215 3689
rect 503530 3680 503536 3732
rect 503588 3720 503594 3732
rect 514113 3723 514171 3729
rect 514113 3720 514125 3723
rect 503588 3692 514125 3720
rect 503588 3680 503594 3692
rect 514113 3689 514125 3692
rect 514159 3689 514171 3723
rect 515600 3720 515628 3760
rect 515677 3757 515689 3791
rect 515723 3788 515735 3791
rect 560846 3788 560852 3800
rect 515723 3760 560852 3788
rect 515723 3757 515735 3760
rect 515677 3751 515735 3757
rect 560846 3748 560852 3760
rect 560904 3748 560910 3800
rect 564434 3720 564440 3732
rect 515600 3692 564440 3720
rect 514113 3683 514171 3689
rect 564434 3680 564440 3692
rect 564492 3680 564498 3732
rect 369452 3624 452700 3652
rect 452749 3655 452807 3661
rect 369452 3612 369458 3624
rect 452749 3621 452761 3655
rect 452795 3652 452807 3655
rect 452795 3624 455460 3652
rect 452795 3621 452807 3624
rect 452749 3615 452807 3621
rect 234672 3556 258074 3584
rect 234672 3544 234678 3556
rect 258258 3544 258264 3596
rect 258316 3584 258322 3596
rect 259270 3584 259276 3596
rect 258316 3556 259276 3584
rect 258316 3544 258322 3556
rect 259270 3544 259276 3556
rect 259328 3544 259334 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 260650 3584 260656 3596
rect 259512 3556 260656 3584
rect 259512 3544 259518 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 261754 3544 261760 3596
rect 261812 3584 261818 3596
rect 262858 3584 262864 3596
rect 261812 3556 262864 3584
rect 261812 3544 261818 3556
rect 262858 3544 262864 3556
rect 262916 3544 262922 3596
rect 273622 3544 273628 3596
rect 273680 3584 273686 3596
rect 274358 3584 274364 3596
rect 273680 3556 274364 3584
rect 273680 3544 273686 3556
rect 274358 3544 274364 3556
rect 274416 3544 274422 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 277213 3587 277271 3593
rect 277213 3553 277225 3587
rect 277259 3584 277271 3587
rect 278038 3584 278044 3596
rect 277259 3556 278044 3584
rect 277259 3553 277271 3556
rect 277213 3547 277271 3553
rect 278038 3544 278044 3556
rect 278096 3544 278102 3596
rect 280706 3544 280712 3596
rect 280764 3584 280770 3596
rect 318150 3584 318156 3596
rect 280764 3556 318156 3584
rect 280764 3544 280770 3556
rect 318150 3544 318156 3556
rect 318208 3544 318214 3596
rect 333882 3544 333888 3596
rect 333940 3584 333946 3596
rect 334710 3584 334716 3596
rect 333940 3556 334716 3584
rect 333940 3544 333946 3556
rect 334710 3544 334716 3556
rect 334768 3544 334774 3596
rect 340874 3544 340880 3596
rect 340932 3584 340938 3596
rect 342162 3584 342168 3596
rect 340932 3556 342168 3584
rect 340932 3544 340938 3556
rect 342162 3544 342168 3556
rect 342220 3544 342226 3596
rect 351638 3544 351644 3596
rect 351696 3584 351702 3596
rect 452473 3587 452531 3593
rect 452473 3584 452485 3587
rect 351696 3556 452485 3584
rect 351696 3544 351702 3556
rect 452473 3553 452485 3556
rect 452519 3553 452531 3587
rect 452473 3547 452531 3553
rect 452841 3587 452899 3593
rect 452841 3553 452853 3587
rect 452887 3584 452899 3587
rect 454405 3587 454463 3593
rect 454405 3584 454417 3587
rect 452887 3556 454417 3584
rect 452887 3553 452899 3556
rect 452841 3547 452899 3553
rect 454405 3553 454417 3556
rect 454451 3553 454463 3587
rect 454405 3547 454463 3553
rect 454494 3544 454500 3596
rect 454552 3584 454558 3596
rect 455322 3584 455328 3596
rect 454552 3556 455328 3584
rect 454552 3544 454558 3556
rect 455322 3544 455328 3556
rect 455380 3544 455386 3596
rect 455432 3584 455460 3624
rect 458082 3612 458088 3664
rect 458140 3652 458146 3664
rect 484578 3652 484584 3664
rect 458140 3624 484584 3652
rect 458140 3612 458146 3624
rect 484578 3612 484584 3624
rect 484636 3612 484642 3664
rect 498010 3612 498016 3664
rect 498068 3652 498074 3664
rect 507670 3652 507676 3664
rect 498068 3624 507676 3652
rect 498068 3612 498074 3624
rect 507670 3612 507676 3624
rect 507728 3612 507734 3664
rect 514662 3612 514668 3664
rect 514720 3652 514726 3664
rect 568022 3652 568028 3664
rect 514720 3624 568028 3652
rect 514720 3612 514726 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 462498 3584 462504 3596
rect 455432 3556 462504 3584
rect 462498 3544 462504 3556
rect 462556 3544 462562 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 510062 3584 510068 3596
rect 467156 3556 510068 3584
rect 467156 3544 467162 3556
rect 510062 3544 510068 3556
rect 510120 3544 510126 3596
rect 510522 3544 510528 3596
rect 510580 3584 510586 3596
rect 515769 3587 515827 3593
rect 515769 3584 515781 3587
rect 510580 3556 515781 3584
rect 510580 3544 510586 3556
rect 515769 3553 515781 3556
rect 515815 3553 515827 3587
rect 571518 3584 571524 3596
rect 515769 3547 515827 3553
rect 515876 3556 571524 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 137278 3516 137284 3528
rect 135312 3488 137284 3516
rect 135312 3476 135318 3488
rect 137278 3476 137284 3488
rect 137336 3476 137342 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144638 3516 144644 3528
rect 143592 3488 144644 3516
rect 143592 3476 143598 3488
rect 144638 3476 144644 3488
rect 144696 3476 144702 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151722 3516 151728 3528
rect 150676 3488 151728 3516
rect 150676 3476 150682 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 155402 3476 155408 3528
rect 155460 3516 155466 3528
rect 155862 3516 155868 3528
rect 155460 3488 155868 3516
rect 155460 3476 155466 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 407390 3516 407396 3528
rect 160204 3488 407396 3516
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 132402 3448 132408 3460
rect 131816 3420 132408 3448
rect 131816 3408 131822 3420
rect 132402 3408 132408 3420
rect 132460 3408 132466 3460
rect 156598 3340 156604 3392
rect 156656 3380 156662 3392
rect 160204 3380 160232 3488
rect 407390 3476 407396 3488
rect 407448 3476 407454 3528
rect 411898 3476 411904 3528
rect 411956 3516 411962 3528
rect 411956 3488 470594 3516
rect 411956 3476 411962 3488
rect 405734 3448 405740 3460
rect 156656 3352 160232 3380
rect 161446 3420 405740 3448
rect 156656 3340 156662 3352
rect 149514 3272 149520 3324
rect 149572 3312 149578 3324
rect 161446 3312 161474 3420
rect 405734 3408 405740 3420
rect 405792 3408 405798 3460
rect 408402 3408 408408 3460
rect 408460 3448 408466 3460
rect 461489 3451 461547 3457
rect 461489 3448 461501 3451
rect 408460 3420 461501 3448
rect 408460 3408 408466 3420
rect 461489 3417 461501 3420
rect 461535 3417 461547 3451
rect 461489 3411 461547 3417
rect 461578 3408 461584 3460
rect 461636 3448 461642 3460
rect 462222 3448 462228 3460
rect 461636 3420 462228 3448
rect 461636 3408 461642 3420
rect 462222 3408 462228 3420
rect 462280 3408 462286 3460
rect 465166 3408 465172 3460
rect 465224 3448 465230 3460
rect 466362 3448 466368 3460
rect 465224 3420 466368 3448
rect 465224 3408 465230 3420
rect 466362 3408 466368 3420
rect 466420 3408 466426 3460
rect 468662 3408 468668 3460
rect 468720 3448 468726 3460
rect 469122 3448 469128 3460
rect 468720 3420 469128 3448
rect 468720 3408 468726 3420
rect 469122 3408 469128 3420
rect 469180 3408 469186 3460
rect 470566 3448 470594 3488
rect 472250 3476 472256 3528
rect 472308 3516 472314 3528
rect 473262 3516 473268 3528
rect 472308 3488 473268 3516
rect 472308 3476 472314 3488
rect 473262 3476 473268 3488
rect 473320 3476 473326 3528
rect 479334 3476 479340 3528
rect 479392 3516 479398 3528
rect 480162 3516 480168 3528
rect 479392 3488 480168 3516
rect 479392 3476 479398 3488
rect 480162 3476 480168 3488
rect 480220 3476 480226 3528
rect 486418 3476 486424 3528
rect 486476 3516 486482 3528
rect 487062 3516 487068 3528
rect 486476 3488 487068 3516
rect 486476 3476 486482 3488
rect 487062 3476 487068 3488
rect 487120 3476 487126 3528
rect 487157 3519 487215 3525
rect 487157 3485 487169 3519
rect 487203 3516 487215 3519
rect 487203 3488 493272 3516
rect 487203 3485 487215 3488
rect 487157 3479 487215 3485
rect 473538 3448 473544 3460
rect 470566 3420 473544 3448
rect 473538 3408 473544 3420
rect 473596 3408 473602 3460
rect 486510 3408 486516 3460
rect 486568 3448 486574 3460
rect 492306 3448 492312 3460
rect 486568 3420 492312 3448
rect 486568 3408 486574 3420
rect 492306 3408 492312 3420
rect 492364 3408 492370 3460
rect 163682 3340 163688 3392
rect 163740 3380 163746 3392
rect 164142 3380 164148 3392
rect 163740 3352 164148 3380
rect 163740 3340 163746 3352
rect 164142 3340 164148 3352
rect 164200 3340 164206 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186222 3380 186228 3392
rect 184992 3352 186228 3380
rect 184992 3340 184998 3352
rect 186222 3340 186228 3352
rect 186280 3340 186286 3392
rect 188522 3340 188528 3392
rect 188580 3380 188586 3392
rect 188982 3380 188988 3392
rect 188580 3352 188988 3380
rect 188580 3340 188586 3352
rect 188982 3340 188988 3352
rect 189040 3340 189046 3392
rect 191098 3340 191104 3392
rect 191156 3380 191162 3392
rect 193214 3380 193220 3392
rect 191156 3352 193220 3380
rect 191156 3340 191162 3352
rect 193214 3340 193220 3352
rect 193272 3340 193278 3392
rect 199102 3340 199108 3392
rect 199160 3380 199166 3392
rect 199930 3380 199936 3392
rect 199160 3352 199936 3380
rect 199160 3340 199166 3352
rect 199930 3340 199936 3352
rect 199988 3340 199994 3392
rect 206186 3340 206192 3392
rect 206244 3380 206250 3392
rect 206830 3380 206836 3392
rect 206244 3352 206836 3380
rect 206244 3340 206250 3352
rect 206830 3340 206836 3352
rect 206888 3340 206894 3392
rect 209774 3340 209780 3392
rect 209832 3380 209838 3392
rect 211062 3380 211068 3392
rect 209832 3352 211068 3380
rect 209832 3340 209838 3352
rect 211062 3340 211068 3352
rect 211120 3340 211126 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 216858 3340 216864 3392
rect 216916 3380 216922 3392
rect 217962 3380 217968 3392
rect 216916 3352 217968 3380
rect 216916 3340 216922 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 241698 3340 241704 3392
rect 241756 3380 241762 3392
rect 242710 3380 242716 3392
rect 241756 3352 242716 3380
rect 241756 3340 241762 3352
rect 242710 3340 242716 3352
rect 242768 3340 242774 3392
rect 245194 3340 245200 3392
rect 245252 3380 245258 3392
rect 246298 3380 246304 3392
rect 245252 3352 246304 3380
rect 245252 3340 245258 3352
rect 246298 3340 246304 3352
rect 246356 3340 246362 3392
rect 254670 3340 254676 3392
rect 254728 3380 254734 3392
rect 255958 3380 255964 3392
rect 254728 3352 255964 3380
rect 254728 3340 254734 3352
rect 255958 3340 255964 3352
rect 256016 3340 256022 3392
rect 270034 3340 270040 3392
rect 270092 3380 270098 3392
rect 277213 3383 277271 3389
rect 277213 3380 277225 3383
rect 270092 3352 277225 3380
rect 270092 3340 270098 3352
rect 277213 3349 277225 3352
rect 277259 3349 277271 3383
rect 277213 3343 277271 3349
rect 305546 3340 305552 3392
rect 305604 3380 305610 3392
rect 306282 3380 306288 3392
rect 305604 3352 306288 3380
rect 305604 3340 305610 3352
rect 306282 3340 306288 3352
rect 306340 3340 306346 3392
rect 312630 3340 312636 3392
rect 312688 3380 312694 3392
rect 342898 3380 342904 3392
rect 312688 3352 342904 3380
rect 312688 3340 312694 3352
rect 342898 3340 342904 3352
rect 342956 3340 342962 3392
rect 348050 3340 348056 3392
rect 348108 3380 348114 3392
rect 378778 3380 378784 3392
rect 348108 3352 378784 3380
rect 348108 3340 348114 3352
rect 378778 3340 378784 3352
rect 378836 3340 378842 3392
rect 397730 3340 397736 3392
rect 397788 3380 397794 3392
rect 460934 3380 460940 3392
rect 397788 3352 460940 3380
rect 397788 3340 397794 3352
rect 460934 3340 460940 3352
rect 460992 3340 460998 3392
rect 461029 3383 461087 3389
rect 461029 3349 461041 3383
rect 461075 3380 461087 3383
rect 467926 3380 467932 3392
rect 461075 3352 467932 3380
rect 461075 3349 461087 3352
rect 461029 3343 461087 3349
rect 467926 3340 467932 3352
rect 467984 3340 467990 3392
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 491202 3380 491208 3392
rect 489972 3352 491208 3380
rect 489972 3340 489978 3352
rect 491202 3340 491208 3352
rect 491260 3340 491266 3392
rect 493244 3380 493272 3488
rect 493502 3476 493508 3528
rect 493560 3516 493566 3528
rect 493962 3516 493968 3528
rect 493560 3488 493968 3516
rect 493560 3476 493566 3488
rect 493962 3476 493968 3488
rect 494020 3476 494026 3528
rect 504358 3476 504364 3528
rect 504416 3516 504422 3528
rect 505370 3516 505376 3528
rect 504416 3488 505376 3516
rect 504416 3476 504422 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 507118 3476 507124 3528
rect 507176 3516 507182 3528
rect 508866 3516 508872 3528
rect 507176 3488 508872 3516
rect 507176 3476 507182 3488
rect 508866 3476 508872 3488
rect 508924 3476 508930 3528
rect 514570 3476 514576 3528
rect 514628 3516 514634 3528
rect 515876 3516 515904 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 514628 3488 515904 3516
rect 514628 3476 514634 3488
rect 516042 3476 516048 3528
rect 516100 3516 516106 3528
rect 575106 3516 575112 3528
rect 516100 3488 575112 3516
rect 516100 3476 516106 3488
rect 575106 3476 575112 3488
rect 575164 3476 575170 3528
rect 493318 3408 493324 3460
rect 493376 3448 493382 3460
rect 494698 3448 494704 3460
rect 493376 3420 494704 3448
rect 493376 3408 493382 3420
rect 494698 3408 494704 3420
rect 494756 3408 494762 3460
rect 500770 3408 500776 3460
rect 500828 3448 500834 3460
rect 514754 3448 514760 3460
rect 500828 3420 514760 3448
rect 500828 3408 500834 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 517422 3408 517428 3460
rect 517480 3448 517486 3460
rect 578602 3448 578608 3460
rect 517480 3420 578608 3448
rect 517480 3408 517486 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 499390 3380 499396 3392
rect 493244 3352 499396 3380
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 499482 3340 499488 3392
rect 499540 3380 499546 3392
rect 511258 3380 511264 3392
rect 499540 3352 511264 3380
rect 499540 3340 499546 3352
rect 511258 3340 511264 3352
rect 511316 3340 511322 3392
rect 539594 3380 539600 3392
rect 513944 3352 539600 3380
rect 149572 3284 161474 3312
rect 149572 3272 149578 3284
rect 162486 3272 162492 3324
rect 162544 3312 162550 3324
rect 170398 3312 170404 3324
rect 162544 3284 170404 3312
rect 162544 3272 162550 3284
rect 170398 3272 170404 3284
rect 170456 3272 170462 3324
rect 192018 3272 192024 3324
rect 192076 3312 192082 3324
rect 192938 3312 192944 3324
rect 192076 3284 192944 3312
rect 192076 3272 192082 3284
rect 192938 3272 192944 3284
rect 192996 3272 193002 3324
rect 223942 3272 223948 3324
rect 224000 3312 224006 3324
rect 228450 3312 228456 3324
rect 224000 3284 228456 3312
rect 224000 3272 224006 3284
rect 228450 3272 228456 3284
rect 228508 3272 228514 3324
rect 401318 3272 401324 3324
rect 401376 3312 401382 3324
rect 470686 3312 470692 3324
rect 401376 3284 470692 3312
rect 401376 3272 401382 3284
rect 470686 3272 470692 3284
rect 470744 3272 470750 3324
rect 495342 3272 495348 3324
rect 495400 3312 495406 3324
rect 497090 3312 497096 3324
rect 495400 3284 497096 3312
rect 495400 3272 495406 3284
rect 497090 3272 497096 3284
rect 497148 3272 497154 3324
rect 506382 3272 506388 3324
rect 506440 3312 506446 3324
rect 513745 3315 513803 3321
rect 513745 3312 513757 3315
rect 506440 3284 513757 3312
rect 506440 3272 506446 3284
rect 513745 3281 513757 3284
rect 513791 3281 513803 3315
rect 513745 3275 513803 3281
rect 283098 3204 283104 3256
rect 283156 3244 283162 3256
rect 284110 3244 284116 3256
rect 283156 3216 284116 3244
rect 283156 3204 283162 3216
rect 284110 3204 284116 3216
rect 284168 3204 284174 3256
rect 404814 3204 404820 3256
rect 404872 3244 404878 3256
rect 470778 3244 470784 3256
rect 404872 3216 470784 3244
rect 404872 3204 404878 3216
rect 470778 3204 470784 3216
rect 470836 3204 470842 3256
rect 506290 3204 506296 3256
rect 506348 3244 506354 3256
rect 513944 3244 513972 3352
rect 539594 3340 539600 3352
rect 539652 3340 539658 3392
rect 514021 3315 514079 3321
rect 514021 3281 514033 3315
rect 514067 3312 514079 3315
rect 536098 3312 536104 3324
rect 514067 3284 536104 3312
rect 514067 3281 514079 3284
rect 514021 3275 514079 3281
rect 536098 3272 536104 3284
rect 536156 3272 536162 3324
rect 532510 3244 532516 3256
rect 506348 3216 513972 3244
rect 514036 3216 532516 3244
rect 506348 3204 506354 3216
rect 141234 3136 141240 3188
rect 141292 3176 141298 3188
rect 142062 3176 142068 3188
rect 141292 3148 142068 3176
rect 141292 3136 141298 3148
rect 142062 3136 142068 3148
rect 142120 3136 142126 3188
rect 175458 3136 175464 3188
rect 175516 3176 175522 3188
rect 178678 3176 178684 3188
rect 175516 3148 178684 3176
rect 175516 3136 175522 3148
rect 178678 3136 178684 3148
rect 178736 3136 178742 3188
rect 291378 3136 291384 3188
rect 291436 3176 291442 3188
rect 298738 3176 298744 3188
rect 291436 3148 298744 3176
rect 291436 3136 291442 3148
rect 298738 3136 298744 3148
rect 298796 3136 298802 3188
rect 422570 3136 422576 3188
rect 422628 3176 422634 3188
rect 423582 3176 423588 3188
rect 422628 3148 423588 3176
rect 422628 3136 422634 3148
rect 423582 3136 423588 3148
rect 423640 3136 423646 3188
rect 474826 3176 474832 3188
rect 427096 3148 474832 3176
rect 186958 3068 186964 3120
rect 187016 3108 187022 3120
rect 189718 3108 189724 3120
rect 187016 3080 189724 3108
rect 187016 3068 187022 3080
rect 189718 3068 189724 3080
rect 189776 3068 189782 3120
rect 418982 3068 418988 3120
rect 419040 3108 419046 3120
rect 427096 3108 427124 3148
rect 474826 3136 474832 3148
rect 474884 3136 474890 3188
rect 505002 3136 505008 3188
rect 505060 3176 505066 3188
rect 514036 3176 514064 3216
rect 532510 3204 532516 3216
rect 532568 3204 532574 3256
rect 505060 3148 514064 3176
rect 514113 3179 514171 3185
rect 505060 3136 505066 3148
rect 514113 3145 514125 3179
rect 514159 3176 514171 3179
rect 529014 3176 529020 3188
rect 514159 3148 529020 3176
rect 514159 3145 514171 3148
rect 514113 3139 514171 3145
rect 529014 3136 529020 3148
rect 529072 3136 529078 3188
rect 476298 3108 476304 3120
rect 419040 3080 427124 3108
rect 427188 3080 476304 3108
rect 419040 3068 419046 3080
rect 174262 3000 174268 3052
rect 174320 3040 174326 3052
rect 175182 3040 175188 3052
rect 174320 3012 175188 3040
rect 174320 3000 174326 3012
rect 175182 3000 175188 3012
rect 175240 3000 175246 3052
rect 284294 3000 284300 3052
rect 284352 3040 284358 3052
rect 285582 3040 285588 3052
rect 284352 3012 285588 3040
rect 284352 3000 284358 3012
rect 285582 3000 285588 3012
rect 285640 3000 285646 3052
rect 415486 3000 415492 3052
rect 415544 3040 415550 3052
rect 416682 3040 416688 3052
rect 415544 3012 416688 3040
rect 415544 3000 415550 3012
rect 416682 3000 416688 3012
rect 416740 3000 416746 3052
rect 426158 3000 426164 3052
rect 426216 3040 426222 3052
rect 427188 3040 427216 3080
rect 476298 3068 476304 3080
rect 476356 3068 476362 3120
rect 503622 3068 503628 3120
rect 503680 3108 503686 3120
rect 525426 3108 525432 3120
rect 503680 3080 525432 3108
rect 503680 3068 503686 3080
rect 525426 3068 525432 3080
rect 525484 3068 525490 3120
rect 426216 3012 427216 3040
rect 426216 3000 426222 3012
rect 429654 3000 429660 3052
rect 429712 3040 429718 3052
rect 477494 3040 477500 3052
rect 429712 3012 477500 3040
rect 429712 3000 429718 3012
rect 477494 3000 477500 3012
rect 477552 3000 477558 3052
rect 490558 3000 490564 3052
rect 490616 3040 490622 3052
rect 498194 3040 498200 3052
rect 490616 3012 498200 3040
rect 490616 3000 490622 3012
rect 498194 3000 498200 3012
rect 498252 3000 498258 3052
rect 502242 3000 502248 3052
rect 502300 3040 502306 3052
rect 521838 3040 521844 3052
rect 502300 3012 521844 3040
rect 502300 3000 502306 3012
rect 521838 3000 521844 3012
rect 521896 3000 521902 3052
rect 171962 2932 171968 2984
rect 172020 2972 172026 2984
rect 179414 2972 179420 2984
rect 172020 2944 179420 2972
rect 172020 2932 172026 2944
rect 179414 2932 179420 2944
rect 179472 2932 179478 2984
rect 440326 2932 440332 2984
rect 440384 2972 440390 2984
rect 441522 2972 441528 2984
rect 440384 2944 441528 2972
rect 440384 2932 440390 2944
rect 441522 2932 441528 2944
rect 441580 2932 441586 2984
rect 447410 2932 447416 2984
rect 447468 2972 447474 2984
rect 448422 2972 448428 2984
rect 447468 2944 448428 2972
rect 447468 2932 447474 2944
rect 448422 2932 448428 2944
rect 448480 2932 448486 2984
rect 478966 2972 478972 2984
rect 448532 2944 478972 2972
rect 436738 2864 436744 2916
rect 436796 2904 436802 2916
rect 448532 2904 448560 2944
rect 478966 2932 478972 2944
rect 479024 2932 479030 2984
rect 500862 2932 500868 2984
rect 500920 2972 500926 2984
rect 518342 2972 518348 2984
rect 500920 2944 518348 2972
rect 500920 2932 500926 2944
rect 518342 2932 518348 2944
rect 518400 2932 518406 2984
rect 481818 2904 481824 2916
rect 436796 2876 448560 2904
rect 448624 2876 481824 2904
rect 436796 2864 436802 2876
rect 443822 2796 443828 2848
rect 443880 2836 443886 2848
rect 448624 2836 448652 2876
rect 481818 2864 481824 2876
rect 481876 2864 481882 2916
rect 443880 2808 448652 2836
rect 443880 2796 443886 2808
rect 450906 2796 450912 2848
rect 450964 2836 450970 2848
rect 483014 2836 483020 2848
rect 450964 2808 483020 2836
rect 450964 2796 450970 2808
rect 483014 2796 483020 2808
rect 483072 2796 483078 2848
<< via1 >>
rect 430488 700408 430540 700460
rect 462320 700408 462372 700460
rect 482928 700408 482980 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 393228 700340 393280 700392
rect 413652 700340 413704 700392
rect 444288 700340 444340 700392
rect 478512 700340 478564 700392
rect 495348 700340 495400 700392
rect 543464 700340 543516 700392
rect 340788 700272 340840 700324
rect 348792 700272 348844 700324
rect 354588 700272 354640 700324
rect 364984 700272 365036 700324
rect 379428 700272 379480 700324
rect 397460 700272 397512 700324
rect 405648 700272 405700 700324
rect 429844 700272 429896 700324
rect 456708 700272 456760 700324
rect 494796 700272 494848 700324
rect 507768 700272 507820 700324
rect 559656 700272 559708 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 328368 699660 328420 699712
rect 332508 699660 332560 699712
rect 522304 696940 522356 696992
rect 580172 696940 580224 696992
rect 522396 683136 522448 683188
rect 580172 683136 580224 683188
rect 522488 670692 522540 670744
rect 580172 670692 580224 670744
rect 300768 655460 300820 655512
rect 302332 655460 302384 655512
rect 353576 655460 353628 655512
rect 354588 655460 354640 655512
rect 443184 655460 443236 655512
rect 444288 655460 444340 655512
rect 455972 655460 456024 655512
rect 456708 655460 456760 655512
rect 481640 655460 481692 655512
rect 482928 655460 482980 655512
rect 494428 654984 494480 655036
rect 495348 654984 495400 655036
rect 41328 654916 41380 654968
rect 97540 654916 97592 654968
rect 106188 654916 106240 654968
rect 148784 654916 148836 654968
rect 171048 654916 171100 654968
rect 199936 654916 199988 654968
rect 24768 654848 24820 654900
rect 84752 654848 84804 654900
rect 89628 654848 89680 654900
rect 135996 654848 136048 654900
rect 154488 654848 154540 654900
rect 187148 654848 187200 654900
rect 219348 654848 219400 654900
rect 238300 654848 238352 654900
rect 8208 654780 8260 654832
rect 72976 654780 73028 654832
rect 73068 654780 73120 654832
rect 123116 654780 123168 654832
rect 137928 654780 137980 654832
rect 174360 654780 174412 654832
rect 202788 654780 202840 654832
rect 225512 654780 225564 654832
rect 235908 654780 235960 654832
rect 251180 654780 251232 654832
rect 267648 654780 267700 654832
rect 276756 654780 276808 654832
rect 404820 654780 404872 654832
rect 405648 654780 405700 654832
rect 392032 654576 392084 654628
rect 393228 654576 393280 654628
rect 284208 654372 284260 654424
rect 289544 654372 289596 654424
rect 507216 654372 507268 654424
rect 507768 654372 507820 654424
rect 522304 643084 522356 643136
rect 580172 643084 580224 643136
rect 3424 641656 3476 641708
rect 69020 641656 69072 641708
rect 522396 630640 522448 630692
rect 580172 630640 580224 630692
rect 3516 630572 3568 630624
rect 69020 630572 69072 630624
rect 3608 619556 3660 619608
rect 69020 619556 69072 619608
rect 522488 616836 522540 616888
rect 580172 616836 580224 616888
rect 3424 597456 3476 597508
rect 69020 597456 69072 597508
rect 522304 590656 522356 590708
rect 579804 590656 579856 590708
rect 3516 585080 3568 585132
rect 69020 585080 69072 585132
rect 522396 576852 522448 576904
rect 580172 576852 580224 576904
rect 3608 573996 3660 574048
rect 69020 573996 69072 574048
rect 522488 563048 522540 563100
rect 579804 563048 579856 563100
rect 3424 551964 3476 552016
rect 69020 551964 69072 552016
rect 3516 540880 3568 540932
rect 69020 540880 69072 540932
rect 522304 536800 522356 536852
rect 580172 536800 580224 536852
rect 3608 529864 3660 529916
rect 69020 529864 69072 529916
rect 522396 524424 522448 524476
rect 580172 524424 580224 524476
rect 522304 510620 522356 510672
rect 580172 510620 580224 510672
rect 3424 507764 3476 507816
rect 69020 507764 69072 507816
rect 3516 496748 3568 496800
rect 69020 496748 69072 496800
rect 3424 485732 3476 485784
rect 69020 485732 69072 485784
rect 522304 484372 522356 484424
rect 580172 484372 580224 484424
rect 522396 470568 522448 470620
rect 579988 470568 580040 470620
rect 3424 462272 3476 462324
rect 69020 462272 69072 462324
rect 522304 456764 522356 456816
rect 580172 456764 580224 456816
rect 3516 451188 3568 451240
rect 69020 451188 69072 451240
rect 3424 440172 3476 440224
rect 69020 440172 69072 440224
rect 522948 430584 523000 430636
rect 580172 430584 580224 430636
rect 522948 418140 523000 418192
rect 580172 418140 580224 418192
rect 3332 418072 3384 418124
rect 69020 418072 69072 418124
rect 3424 407056 3476 407108
rect 69020 407056 69072 407108
rect 522028 404336 522080 404388
rect 580172 404336 580224 404388
rect 2872 395972 2924 396024
rect 69020 395972 69072 396024
rect 522948 378768 523000 378820
rect 580172 378768 580224 378820
rect 3424 372580 3476 372632
rect 69020 372580 69072 372632
rect 522948 365644 523000 365696
rect 580172 365644 580224 365696
rect 3424 361564 3476 361616
rect 69020 361564 69072 361616
rect 522948 353200 523000 353252
rect 580172 353200 580224 353252
rect 2872 349120 2924 349172
rect 69020 349120 69072 349172
rect 2872 327088 2924 327140
rect 69020 327088 69072 327140
rect 522304 325592 522356 325644
rect 580172 325592 580224 325644
rect 3516 316004 3568 316056
rect 69020 316004 69072 316056
rect 522304 313216 522356 313268
rect 580172 313216 580224 313268
rect 3424 304988 3476 305040
rect 69020 304988 69072 305040
rect 522304 299412 522356 299464
rect 580172 299412 580224 299464
rect 3424 282888 3476 282940
rect 69020 282888 69072 282940
rect 522396 273164 522448 273216
rect 580172 273164 580224 273216
rect 3516 271872 3568 271924
rect 69020 271872 69072 271924
rect 3424 260856 3476 260908
rect 69020 260856 69072 260908
rect 522304 259360 522356 259412
rect 580172 259360 580224 259412
rect 522396 245556 522448 245608
rect 580172 245556 580224 245608
rect 3516 238756 3568 238808
rect 69020 238756 69072 238808
rect 522304 233180 522356 233232
rect 579988 233180 580040 233232
rect 3608 226312 3660 226364
rect 69020 226312 69072 226364
rect 522396 219376 522448 219428
rect 580172 219376 580224 219428
rect 3424 215296 3476 215348
rect 69020 215296 69072 215348
rect 522304 206932 522356 206984
rect 579804 206932 579856 206984
rect 3608 193196 3660 193248
rect 69020 193196 69072 193248
rect 522488 193128 522540 193180
rect 580172 193128 580224 193180
rect 3516 182180 3568 182232
rect 69020 182180 69072 182232
rect 522396 179324 522448 179376
rect 580172 179324 580224 179376
rect 3424 171096 3476 171148
rect 69020 171096 69072 171148
rect 522304 166948 522356 167000
rect 580172 166948 580224 167000
rect 522488 153144 522540 153196
rect 580172 153144 580224 153196
rect 3700 149064 3752 149116
rect 69020 149064 69072 149116
rect 522396 139340 522448 139392
rect 580172 139340 580224 139392
rect 3608 137980 3660 138032
rect 69020 137980 69072 138032
rect 3516 126964 3568 127016
rect 69020 126964 69072 127016
rect 522304 126896 522356 126948
rect 580172 126896 580224 126948
rect 3424 114520 3476 114572
rect 69020 114520 69072 114572
rect 522580 113092 522632 113144
rect 579804 113092 579856 113144
rect 3792 103504 3844 103556
rect 69020 103504 69072 103556
rect 522488 100648 522540 100700
rect 580172 100648 580224 100700
rect 3700 92488 3752 92540
rect 69020 92488 69072 92540
rect 522396 86912 522448 86964
rect 580172 86912 580224 86964
rect 3608 81404 3660 81456
rect 69020 81404 69072 81456
rect 522304 73108 522356 73160
rect 580172 73108 580224 73160
rect 3516 70388 3568 70440
rect 69020 70388 69072 70440
rect 3424 60732 3476 60784
rect 69020 60732 69072 60784
rect 522672 60664 522724 60716
rect 580172 60664 580224 60716
rect 295340 59780 295392 59832
rect 296316 59780 296368 59832
rect 313372 59780 313424 59832
rect 314532 59780 314584 59832
rect 324320 59780 324372 59832
rect 325388 59780 325440 59832
rect 427820 59780 427872 59832
rect 428980 59780 429032 59832
rect 430580 59780 430632 59832
rect 431740 59780 431792 59832
rect 436100 59780 436152 59832
rect 437168 59780 437220 59832
rect 438860 59780 438912 59832
rect 439928 59780 439980 59832
rect 456800 59780 456852 59832
rect 458052 59780 458104 59832
rect 467840 59780 467892 59832
rect 469000 59780 469052 59832
rect 155868 57876 155920 57928
rect 291752 57876 291804 57928
rect 383660 57876 383712 57928
rect 384856 57876 384908 57928
rect 469128 57876 469180 57928
rect 487988 57876 488040 57928
rect 153108 57808 153160 57860
rect 290832 57808 290884 57860
rect 375472 57808 375524 57860
rect 443644 57808 443696 57860
rect 473268 57808 473320 57860
rect 488908 57808 488960 57860
rect 136548 57740 136600 57792
rect 170864 57740 170916 57792
rect 184664 57740 184716 57792
rect 186964 57740 187016 57792
rect 187332 57740 187384 57792
rect 200120 57740 200172 57792
rect 201316 57740 201368 57792
rect 218244 57740 218296 57792
rect 222844 57740 222896 57792
rect 225512 57740 225564 57792
rect 233884 57740 233936 57792
rect 234620 57740 234672 57792
rect 374644 57740 374696 57792
rect 380900 57740 380952 57792
rect 449164 57740 449216 57792
rect 466368 57740 466420 57792
rect 487160 57740 487212 57792
rect 148968 57672 149020 57724
rect 289912 57672 289964 57724
rect 377404 57672 377456 57724
rect 455420 57672 455472 57724
rect 462228 57672 462280 57724
rect 486240 57672 486292 57724
rect 144828 57604 144880 57656
rect 288992 57604 289044 57656
rect 305644 57604 305696 57656
rect 321560 57604 321612 57656
rect 332600 57604 332652 57656
rect 333520 57604 333572 57656
rect 335360 57604 335412 57656
rect 336280 57604 336332 57656
rect 339960 57604 340012 57656
rect 340788 57604 340840 57656
rect 340880 57604 340932 57656
rect 342076 57604 342128 57656
rect 342720 57604 342772 57656
rect 343548 57604 343600 57656
rect 343640 57604 343692 57656
rect 344928 57604 344980 57656
rect 345480 57604 345532 57656
rect 346308 57604 346360 57656
rect 346400 57604 346452 57656
rect 347596 57604 347648 57656
rect 348148 57604 348200 57656
rect 348976 57604 349028 57656
rect 350908 57604 350960 57656
rect 351736 57604 351788 57656
rect 353668 57604 353720 57656
rect 354588 57604 354640 57656
rect 355416 57604 355468 57656
rect 355968 57604 356020 57656
rect 356336 57604 356388 57656
rect 357256 57604 357308 57656
rect 358176 57604 358228 57656
rect 358728 57604 358780 57656
rect 359096 57604 359148 57656
rect 360016 57604 360068 57656
rect 360936 57604 360988 57656
rect 361488 57604 361540 57656
rect 363604 57604 363656 57656
rect 364248 57604 364300 57656
rect 364524 57604 364576 57656
rect 365536 57604 365588 57656
rect 366364 57604 366416 57656
rect 367008 57604 367060 57656
rect 367284 57604 367336 57656
rect 368388 57604 368440 57656
rect 369032 57604 369084 57656
rect 369768 57604 369820 57656
rect 369952 57604 370004 57656
rect 371056 57604 371108 57656
rect 371792 57604 371844 57656
rect 372528 57604 372580 57656
rect 372712 57604 372764 57656
rect 373816 57604 373868 57656
rect 374552 57604 374604 57656
rect 375288 57604 375340 57656
rect 377220 57604 377272 57656
rect 378048 57604 378100 57656
rect 378140 57604 378192 57656
rect 379336 57604 379388 57656
rect 379980 57604 380032 57656
rect 483664 57604 483716 57656
rect 496268 57604 496320 57656
rect 497464 57604 497516 57656
rect 499028 57604 499080 57656
rect 499488 57604 499540 57656
rect 499948 57604 500000 57656
rect 500776 57604 500828 57656
rect 502616 57604 502668 57656
rect 503628 57604 503680 57656
rect 505376 57604 505428 57656
rect 506388 57604 506440 57656
rect 508136 57604 508188 57656
rect 509056 57604 509108 57656
rect 509884 57604 509936 57656
rect 510528 57604 510580 57656
rect 510804 57604 510856 57656
rect 511816 57604 511868 57656
rect 512644 57604 512696 57656
rect 513288 57604 513340 57656
rect 513564 57604 513616 57656
rect 514668 57604 514720 57656
rect 515404 57604 515456 57656
rect 516048 57604 516100 57656
rect 142068 57536 142120 57588
rect 288164 57536 288216 57588
rect 288256 57536 288308 57588
rect 300860 57536 300912 57588
rect 320824 57536 320876 57588
rect 444380 57536 444432 57588
rect 449900 57536 449952 57588
rect 450728 57536 450780 57588
rect 452660 57536 452712 57588
rect 453488 57536 453540 57588
rect 455328 57536 455380 57588
rect 484400 57536 484452 57588
rect 497188 57536 497240 57588
rect 498108 57536 498160 57588
rect 516232 57536 516284 57588
rect 517428 57536 517480 57588
rect 140688 57468 140740 57520
rect 171784 57468 171836 57520
rect 183744 57468 183796 57520
rect 184848 57468 184900 57520
rect 186412 57468 186464 57520
rect 187608 57468 187660 57520
rect 133788 57400 133840 57452
rect 170036 57400 170088 57452
rect 188252 57400 188304 57452
rect 191012 57468 191064 57520
rect 191748 57468 191800 57520
rect 191932 57468 191984 57520
rect 193036 57468 193088 57520
rect 193680 57468 193732 57520
rect 194508 57468 194560 57520
rect 194600 57468 194652 57520
rect 195888 57468 195940 57520
rect 196440 57468 196492 57520
rect 197268 57468 197320 57520
rect 197360 57468 197412 57520
rect 198648 57468 198700 57520
rect 199200 57468 199252 57520
rect 200028 57468 200080 57520
rect 200948 57468 201000 57520
rect 201408 57468 201460 57520
rect 201868 57468 201920 57520
rect 202788 57468 202840 57520
rect 203708 57468 203760 57520
rect 204168 57468 204220 57520
rect 204628 57468 204680 57520
rect 205548 57468 205600 57520
rect 206468 57468 206520 57520
rect 206928 57468 206980 57520
rect 209136 57468 209188 57520
rect 209688 57468 209740 57520
rect 212816 57468 212868 57520
rect 213736 57468 213788 57520
rect 214656 57468 214708 57520
rect 215208 57468 215260 57520
rect 215484 57468 215536 57520
rect 216496 57468 216548 57520
rect 217324 57468 217376 57520
rect 217968 57468 218020 57520
rect 200120 57400 200172 57452
rect 211896 57400 211948 57452
rect 219992 57468 220044 57520
rect 220084 57468 220136 57520
rect 220728 57468 220780 57520
rect 222752 57468 222804 57520
rect 223396 57468 223448 57520
rect 223672 57468 223724 57520
rect 224868 57468 224920 57520
rect 229192 57468 229244 57520
rect 230296 57468 230348 57520
rect 230940 57468 230992 57520
rect 231768 57468 231820 57520
rect 231860 57468 231912 57520
rect 233056 57468 233108 57520
rect 233700 57468 233752 57520
rect 234528 57468 234580 57520
rect 237288 57468 237340 57520
rect 238024 57468 238076 57520
rect 219164 57400 219216 57452
rect 221924 57400 221976 57452
rect 231124 57400 231176 57452
rect 236460 57400 236512 57452
rect 384488 57468 384540 57520
rect 384948 57468 385000 57520
rect 385408 57468 385460 57520
rect 386328 57468 386380 57520
rect 387248 57468 387300 57520
rect 387708 57468 387760 57520
rect 388168 57468 388220 57520
rect 388996 57468 389048 57520
rect 390008 57468 390060 57520
rect 390468 57468 390520 57520
rect 390928 57468 390980 57520
rect 391756 57468 391808 57520
rect 392676 57468 392728 57520
rect 393228 57468 393280 57520
rect 393596 57468 393648 57520
rect 394516 57468 394568 57520
rect 395436 57468 395488 57520
rect 395988 57468 396040 57520
rect 396356 57468 396408 57520
rect 397368 57468 397420 57520
rect 398196 57468 398248 57520
rect 398748 57468 398800 57520
rect 399024 57468 399076 57520
rect 400128 57468 400180 57520
rect 238208 57400 238260 57452
rect 238668 57400 238720 57452
rect 240048 57400 240100 57452
rect 240784 57400 240836 57452
rect 240968 57400 241020 57452
rect 241428 57400 241480 57452
rect 241888 57400 241940 57452
rect 242716 57400 242768 57452
rect 243728 57400 243780 57452
rect 244188 57400 244240 57452
rect 244556 57400 244608 57452
rect 245568 57400 245620 57452
rect 246396 57400 246448 57452
rect 246948 57400 247000 57452
rect 247316 57400 247368 57452
rect 248236 57400 248288 57452
rect 394792 57400 394844 57452
rect 404452 57468 404504 57520
rect 412732 57468 412784 57520
rect 413468 57468 413520 57520
rect 415400 57468 415452 57520
rect 416228 57468 416280 57520
rect 418160 57468 418212 57520
rect 418988 57468 419040 57520
rect 435364 57468 435416 57520
rect 440792 57468 440844 57520
rect 448428 57468 448480 57520
rect 482560 57468 482612 57520
rect 403624 57400 403676 57452
rect 438032 57400 438084 57452
rect 441528 57400 441580 57452
rect 480720 57400 480772 57452
rect 487068 57400 487120 57452
rect 492680 57400 492732 57452
rect 501696 57400 501748 57452
rect 502248 57400 502300 57452
rect 504456 57400 504508 57452
rect 505008 57400 505060 57452
rect 507216 57400 507268 57452
rect 507768 57400 507820 57452
rect 2688 57332 2740 57384
rect 72792 57332 72844 57384
rect 129648 57332 129700 57384
rect 169116 57332 169168 57384
rect 188344 57332 188396 57384
rect 408960 57332 409012 57384
rect 421564 57332 421616 57384
rect 427176 57332 427228 57384
rect 433248 57332 433300 57384
rect 478880 57332 478932 57384
rect 480168 57332 480220 57384
rect 490748 57332 490800 57384
rect 126888 57264 126940 57316
rect 168196 57264 168248 57316
rect 173164 57264 173216 57316
rect 407120 57264 407172 57316
rect 423588 57264 423640 57316
rect 476212 57264 476264 57316
rect 482928 57264 482980 57316
rect 491668 57332 491720 57384
rect 491208 57264 491260 57316
rect 493508 57264 493560 57316
rect 1308 57196 1360 57248
rect 72976 57196 73028 57248
rect 162124 57196 162176 57248
rect 405372 57196 405424 57248
rect 416688 57196 416740 57248
rect 474372 57196 474424 57248
rect 476028 57196 476080 57248
rect 489920 57196 489972 57248
rect 169024 57128 169076 57180
rect 287244 57128 287296 57180
rect 382740 57128 382792 57180
rect 383568 57128 383620 57180
rect 389824 57128 389876 57180
rect 400864 57128 400916 57180
rect 144736 57060 144788 57112
rect 172704 57060 172756 57112
rect 189172 57060 189224 57112
rect 190276 57060 190328 57112
rect 196624 57060 196676 57112
rect 210976 57060 211028 57112
rect 151728 56992 151780 57044
rect 174544 56992 174596 57044
rect 207388 56992 207440 57044
rect 208216 56992 208268 57044
rect 210056 56992 210108 57044
rect 214564 56992 214616 57044
rect 228364 56992 228416 57044
rect 239128 56992 239180 57044
rect 249156 56992 249208 57044
rect 249708 56992 249760 57044
rect 250076 56992 250128 57044
rect 250996 56992 251048 57044
rect 251824 56992 251876 57044
rect 252468 56992 252520 57044
rect 252744 56992 252796 57044
rect 253848 56992 253900 57044
rect 254584 56992 254636 57044
rect 255228 56992 255280 57044
rect 255504 56992 255556 57044
rect 256516 56992 256568 57044
rect 257344 56992 257396 57044
rect 257988 56992 258040 57044
rect 258264 57060 258316 57112
rect 259368 57060 259420 57112
rect 260012 57060 260064 57112
rect 260748 57060 260800 57112
rect 262772 57060 262824 57112
rect 263508 57060 263560 57112
rect 263692 57060 263744 57112
rect 264888 57060 264940 57112
rect 266360 57060 266412 57112
rect 267556 57060 267608 57112
rect 268200 57060 268252 57112
rect 269028 57060 269080 57112
rect 269120 57060 269172 57112
rect 270316 57060 270368 57112
rect 270960 57060 271012 57112
rect 271788 57060 271840 57112
rect 271880 57060 271932 57112
rect 273168 57060 273220 57112
rect 273628 57060 273680 57112
rect 274548 57060 274600 57112
rect 275468 57060 275520 57112
rect 275928 57060 275980 57112
rect 276388 57060 276440 57112
rect 277308 57060 277360 57112
rect 278228 57060 278280 57112
rect 278688 57060 278740 57112
rect 279148 57060 279200 57112
rect 279976 57060 280028 57112
rect 280988 57060 281040 57112
rect 281448 57060 281500 57112
rect 281816 57060 281868 57112
rect 282828 57060 282880 57112
rect 283656 57060 283708 57112
rect 284208 57060 284260 57112
rect 286324 57060 286376 57112
rect 319904 57060 319956 57112
rect 264244 56992 264296 57044
rect 147588 56924 147640 56976
rect 173624 56924 173676 56976
rect 259092 56924 259144 56976
rect 287796 56992 287848 57044
rect 288440 56992 288492 57044
rect 292672 56992 292724 57044
rect 264612 56924 264664 56976
rect 291936 56924 291988 56976
rect 158628 56856 158680 56908
rect 176384 56856 176436 56908
rect 228272 56856 228324 56908
rect 229008 56856 229060 56908
rect 161388 56788 161440 56840
rect 177304 56788 177356 56840
rect 165528 56720 165580 56772
rect 178132 56720 178184 56772
rect 260932 56720 260984 56772
rect 289084 56856 289136 56908
rect 309232 56720 309284 56772
rect 309968 56720 310020 56772
rect 347228 56720 347280 56772
rect 347688 56720 347740 56772
rect 349988 56720 350040 56772
rect 350448 56720 350500 56772
rect 352748 56720 352800 56772
rect 353208 56720 353260 56772
rect 361764 56720 361816 56772
rect 362776 56720 362828 56772
rect 166264 56652 166316 56704
rect 175464 56652 175516 56704
rect 178684 56652 178736 56704
rect 180892 56652 180944 56704
rect 185584 56652 185636 56704
rect 191104 56652 191156 56704
rect 180064 56584 180116 56636
rect 181812 56584 181864 56636
rect 221004 56584 221056 56636
rect 287704 56584 287756 56636
rect 288256 56584 288308 56636
rect 291844 56584 291896 56636
rect 297180 56584 297232 56636
rect 429844 56584 429896 56636
rect 434444 56584 434496 56636
rect 262864 56312 262916 56364
rect 318984 56312 319036 56364
rect 382924 56312 382976 56364
rect 456248 56312 456300 56364
rect 331220 56244 331272 56296
rect 363604 56244 363656 56296
rect 451648 56244 451700 56296
rect 177304 56176 177356 56228
rect 294512 56176 294564 56228
rect 322204 56176 322256 56228
rect 441712 56176 441764 56228
rect 170404 56108 170456 56160
rect 293592 56108 293644 56160
rect 318064 56108 318116 56160
rect 445300 56108 445352 56160
rect 447140 56108 447192 56160
rect 448060 56108 448112 56160
rect 280804 56040 280856 56092
rect 433524 56040 433576 56092
rect 261852 55972 261904 56024
rect 489184 55972 489236 56024
rect 265532 55904 265584 55956
rect 504364 55904 504416 55956
rect 137284 55836 137336 55888
rect 402612 55836 402664 55888
rect 298100 55700 298152 55752
rect 299020 55700 299072 55752
rect 226432 54612 226484 54664
rect 351920 54612 351972 54664
rect 160008 54544 160060 54596
rect 288440 54544 288492 54596
rect 340144 54544 340196 54596
rect 447232 54544 447284 54596
rect 143448 54476 143500 54528
rect 394792 54476 394844 54528
rect 233884 50328 233936 50380
rect 349160 50328 349212 50380
rect 522580 46860 522632 46912
rect 580172 46860 580224 46912
rect 376024 40672 376076 40724
rect 454040 40672 454092 40724
rect 371884 39312 371936 39364
rect 452752 39312 452804 39364
rect 260104 37884 260156 37936
rect 427912 37884 427964 37936
rect 342904 36524 342956 36576
rect 447140 36524 447192 36576
rect 184204 35164 184256 35216
rect 298192 35164 298244 35216
rect 298744 35164 298796 35216
rect 441620 35164 441672 35216
rect 246304 33736 246356 33788
rect 430672 33736 430724 33788
rect 522488 33056 522540 33108
rect 580172 33056 580224 33108
rect 227536 32376 227588 32428
rect 425152 32376 425204 32428
rect 240784 31016 240836 31068
rect 405832 31016 405884 31068
rect 294604 29588 294656 29640
rect 438952 29588 439004 29640
rect 142804 28228 142856 28280
rect 402980 28228 403032 28280
rect 271144 26868 271196 26920
rect 431960 26868 432012 26920
rect 169668 25508 169720 25560
rect 295432 25508 295484 25560
rect 295984 25508 296036 25560
rect 436192 25508 436244 25560
rect 238024 24080 238076 24132
rect 394700 24080 394752 24132
rect 224776 22720 224828 22772
rect 345020 22720 345072 22772
rect 358084 22720 358136 22772
rect 448520 22720 448572 22772
rect 222844 21428 222896 21480
rect 320180 21428 320232 21480
rect 238024 21360 238076 21412
rect 423680 21360 423732 21412
rect 522396 20612 522448 20664
rect 579988 20612 580040 20664
rect 268936 20000 268988 20052
rect 320272 20000 320324 20052
rect 214564 19932 214616 19984
rect 288440 19932 288492 19984
rect 323584 19932 323636 19984
rect 443000 19932 443052 19984
rect 357256 18708 357308 18760
rect 407212 18708 407264 18760
rect 231124 18640 231176 18692
rect 334072 18640 334124 18692
rect 356704 18640 356756 18692
rect 449992 18640 450044 18692
rect 231676 18572 231728 18624
rect 421564 18572 421616 18624
rect 214564 17484 214616 17536
rect 299480 17484 299532 17536
rect 378784 17416 378836 17468
rect 456892 17416 456944 17468
rect 213736 17348 213788 17400
rect 299480 17348 299532 17400
rect 379336 17348 379388 17400
rect 486424 17348 486476 17400
rect 298836 17280 298888 17332
rect 434720 17280 434772 17332
rect 278044 17212 278096 17264
rect 436100 17212 436152 17264
rect 224224 16124 224276 16176
rect 298100 16124 298152 16176
rect 267004 16056 267056 16108
rect 430580 16056 430632 16108
rect 249064 15988 249116 16040
rect 427820 15988 427872 16040
rect 228456 15920 228508 15972
rect 425060 15920 425112 15972
rect 267556 15852 267608 15904
rect 507124 15852 507176 15904
rect 259276 14900 259328 14952
rect 317420 14900 317472 14952
rect 173808 14832 173860 14884
rect 295340 14832 295392 14884
rect 318156 14832 318208 14884
rect 438860 14832 438912 14884
rect 274364 14764 274416 14816
rect 403624 14764 403676 14816
rect 229008 14696 229060 14748
rect 359464 14696 359516 14748
rect 360844 14696 360896 14748
rect 449900 14696 449952 14748
rect 242716 14628 242768 14680
rect 412640 14628 412692 14680
rect 235908 14560 235960 14612
rect 387800 14560 387852 14612
rect 242716 14492 242768 14544
rect 429200 14492 429252 14544
rect 264888 14424 264940 14476
rect 490564 14424 490616 14476
rect 255964 13676 256016 13728
rect 316132 13676 316184 13728
rect 228364 13608 228416 13660
rect 324412 13608 324464 13660
rect 217968 13540 218020 13592
rect 317328 13540 317380 13592
rect 383568 13540 383620 13592
rect 467104 13540 467156 13592
rect 224868 13472 224920 13524
rect 340880 13472 340932 13524
rect 378048 13472 378100 13524
rect 488816 13472 488868 13524
rect 220728 13404 220780 13456
rect 327080 13404 327132 13456
rect 334716 13404 334768 13456
rect 452660 13404 452712 13456
rect 285588 13336 285640 13388
rect 435364 13336 435416 13388
rect 238668 13268 238720 13320
rect 398932 13268 398984 13320
rect 260656 13200 260708 13252
rect 429844 13200 429896 13252
rect 291936 13132 291988 13184
rect 501328 13132 501380 13184
rect 263508 13064 263560 13116
rect 493324 13064 493376 13116
rect 277124 12384 277176 12436
rect 321652 12384 321704 12436
rect 215208 12316 215260 12368
rect 306380 12316 306432 12368
rect 216496 12248 216548 12300
rect 309784 12248 309836 12300
rect 357348 12248 357400 12300
rect 410800 12248 410852 12300
rect 216588 12180 216640 12232
rect 313832 12180 313884 12232
rect 376668 12180 376720 12232
rect 484492 12180 484544 12232
rect 223488 12112 223540 12164
rect 338672 12112 338724 12164
rect 379428 12112 379480 12164
rect 495440 12112 495492 12164
rect 227628 12044 227680 12096
rect 356336 12044 356388 12096
rect 382188 12044 382240 12096
rect 506480 12044 506532 12096
rect 213828 11976 213880 12028
rect 303160 11976 303212 12028
rect 306288 11976 306340 12028
rect 445760 11976 445812 12028
rect 241428 11908 241480 11960
rect 409144 11908 409196 11960
rect 287796 11840 287848 11892
rect 480536 11840 480588 11892
rect 289084 11772 289136 11824
rect 487160 11772 487212 11824
rect 260748 11704 260800 11756
rect 483664 11704 483716 11756
rect 192944 10956 192996 11008
rect 416780 10956 416832 11008
rect 188988 10888 189040 10940
rect 415400 10888 415452 10940
rect 186228 10820 186280 10872
rect 415492 10820 415544 10872
rect 182088 10752 182140 10804
rect 414020 10752 414072 10804
rect 177856 10684 177908 10736
rect 412732 10684 412784 10736
rect 175188 10616 175240 10668
rect 412824 10616 412876 10668
rect 170772 10548 170824 10600
rect 411260 10548 411312 10600
rect 168288 10480 168340 10532
rect 410064 10480 410116 10532
rect 164148 10412 164200 10464
rect 409972 10412 410024 10464
rect 132408 10344 132460 10396
rect 401600 10344 401652 10396
rect 128176 10276 128228 10328
rect 400220 10276 400272 10328
rect 195612 10208 195664 10260
rect 418252 10208 418304 10260
rect 199936 10140 199988 10192
rect 418160 10140 418212 10192
rect 202604 10072 202656 10124
rect 419540 10072 419592 10124
rect 206836 10004 206888 10056
rect 419632 10004 419684 10056
rect 211068 9936 211120 9988
rect 420920 9936 420972 9988
rect 213828 9868 213880 9920
rect 422300 9868 422352 9920
rect 217968 9800 218020 9852
rect 422392 9800 422444 9852
rect 284116 9732 284168 9784
rect 324504 9732 324556 9784
rect 222752 9596 222804 9648
rect 309324 9596 309376 9648
rect 365628 9596 365680 9648
rect 442632 9596 442684 9648
rect 219256 9528 219308 9580
rect 307760 9528 307812 9580
rect 367008 9528 367060 9580
rect 446220 9528 446272 9580
rect 215668 9460 215720 9512
rect 306564 9460 306616 9512
rect 368388 9460 368440 9512
rect 449808 9596 449860 9648
rect 212172 9392 212224 9444
rect 306472 9392 306524 9444
rect 368296 9392 368348 9444
rect 453304 9528 453356 9580
rect 449164 9460 449216 9512
rect 502984 9460 503036 9512
rect 208584 9324 208636 9376
rect 305000 9324 305052 9376
rect 369768 9324 369820 9376
rect 456892 9324 456944 9376
rect 205088 9256 205140 9308
rect 303712 9256 303764 9308
rect 371056 9256 371108 9308
rect 460388 9256 460440 9308
rect 201500 9188 201552 9240
rect 303620 9188 303672 9240
rect 371148 9188 371200 9240
rect 463976 9188 464028 9240
rect 197912 9120 197964 9172
rect 302332 9120 302384 9172
rect 372528 9120 372580 9172
rect 467472 9120 467524 9172
rect 194416 9052 194468 9104
rect 300952 9052 301004 9104
rect 373816 9052 373868 9104
rect 471060 9052 471112 9104
rect 134156 8984 134208 9036
rect 285680 8984 285732 9036
rect 373908 8984 373960 9036
rect 474556 8984 474608 9036
rect 130568 8916 130620 8968
rect 284392 8916 284444 8968
rect 375288 8916 375340 8968
rect 478144 8916 478196 8968
rect 226340 8848 226392 8900
rect 309232 8848 309284 8900
rect 365536 8848 365588 8900
rect 439136 8848 439188 8900
rect 229836 8780 229888 8832
rect 310520 8780 310572 8832
rect 364248 8780 364300 8832
rect 435548 8780 435600 8832
rect 233424 8712 233476 8764
rect 310612 8712 310664 8764
rect 362868 8712 362920 8764
rect 432052 8712 432104 8764
rect 237012 8644 237064 8696
rect 311900 8644 311952 8696
rect 362776 8644 362828 8696
rect 428464 8644 428516 8696
rect 240508 8576 240560 8628
rect 313464 8576 313516 8628
rect 361488 8576 361540 8628
rect 424968 8576 425020 8628
rect 244096 8508 244148 8560
rect 313372 8508 313424 8560
rect 360108 8508 360160 8560
rect 421380 8508 421432 8560
rect 247592 8440 247644 8492
rect 314660 8440 314712 8492
rect 360016 8440 360068 8492
rect 417884 8440 417936 8492
rect 251180 8372 251232 8424
rect 316040 8372 316092 8424
rect 358728 8372 358780 8424
rect 414296 8372 414348 8424
rect 249708 8236 249760 8288
rect 441252 8236 441304 8288
rect 443644 8236 443696 8288
rect 481732 8236 481784 8288
rect 250996 8168 251048 8220
rect 445024 8168 445076 8220
rect 251088 8100 251140 8152
rect 448612 8100 448664 8152
rect 252468 8032 252520 8084
rect 452108 8032 452160 8084
rect 253848 7964 253900 8016
rect 455696 7964 455748 8016
rect 253756 7896 253808 7948
rect 459192 7896 459244 7948
rect 255228 7828 255280 7880
rect 462780 7828 462832 7880
rect 256516 7760 256568 7812
rect 466276 7760 466328 7812
rect 256608 7692 256660 7744
rect 469864 7692 469916 7744
rect 257988 7624 258040 7676
rect 473452 7624 473504 7676
rect 259368 7556 259420 7608
rect 476948 7556 477000 7608
rect 248328 7488 248380 7540
rect 437940 7488 437992 7540
rect 248236 7420 248288 7472
rect 434444 7420 434496 7472
rect 246948 7352 247000 7404
rect 430856 7352 430908 7404
rect 245476 7284 245528 7336
rect 427268 7284 427320 7336
rect 245568 7216 245620 7268
rect 423772 7216 423824 7268
rect 244188 7148 244240 7200
rect 420184 7148 420236 7200
rect 242808 7080 242860 7132
rect 416412 7080 416464 7132
rect 126980 7012 127032 7064
rect 284300 7012 284352 7064
rect 355968 7012 356020 7064
rect 403624 7012 403676 7064
rect 279516 6808 279568 6860
rect 322940 6808 322992 6860
rect 350448 6808 350500 6860
rect 382372 6808 382424 6860
rect 522304 6808 522356 6860
rect 580172 6808 580224 6860
rect 209688 6740 209740 6792
rect 285404 6740 285456 6792
rect 286600 6740 286652 6792
rect 324320 6740 324372 6792
rect 325608 6740 325660 6792
rect 335452 6740 335504 6792
rect 351736 6740 351788 6792
rect 385960 6740 386012 6792
rect 391848 6740 391900 6792
rect 545488 6740 545540 6792
rect 220084 6672 220136 6724
rect 296076 6672 296128 6724
rect 297272 6672 297324 6724
rect 327264 6672 327316 6724
rect 351828 6672 351880 6724
rect 389456 6672 389508 6724
rect 393228 6672 393280 6724
rect 549076 6672 549128 6724
rect 190828 6604 190880 6656
rect 287704 6604 287756 6656
rect 290188 6604 290240 6656
rect 325700 6604 325752 6656
rect 342168 6604 342220 6656
rect 350448 6604 350500 6656
rect 353208 6604 353260 6656
rect 393044 6604 393096 6656
rect 394516 6604 394568 6656
rect 552664 6604 552716 6656
rect 176660 6536 176712 6588
rect 291844 6536 291896 6588
rect 293684 6536 293736 6588
rect 327172 6536 327224 6588
rect 343548 6536 343600 6588
rect 354036 6536 354088 6588
rect 354588 6536 354640 6588
rect 230296 6468 230348 6520
rect 363512 6468 363564 6520
rect 230388 6400 230440 6452
rect 367008 6400 367060 6452
rect 394608 6536 394660 6588
rect 556160 6536 556212 6588
rect 395896 6468 395948 6520
rect 559748 6468 559800 6520
rect 396540 6400 396592 6452
rect 397368 6400 397420 6452
rect 563244 6400 563296 6452
rect 231768 6332 231820 6384
rect 370596 6332 370648 6384
rect 397276 6332 397328 6384
rect 566832 6332 566884 6384
rect 233056 6264 233108 6316
rect 374092 6264 374144 6316
rect 374644 6264 374696 6316
rect 384764 6264 384816 6316
rect 398748 6264 398800 6316
rect 570328 6264 570380 6316
rect 233148 6196 233200 6248
rect 377680 6196 377732 6248
rect 391756 6196 391808 6248
rect 400128 6196 400180 6248
rect 573916 6196 573968 6248
rect 234528 6128 234580 6180
rect 381176 6128 381228 6180
rect 384856 6128 384908 6180
rect 399944 6128 399996 6180
rect 400036 6128 400088 6180
rect 577412 6128 577464 6180
rect 272432 6060 272484 6112
rect 305644 6060 305696 6112
rect 307944 6060 307996 6112
rect 329932 6060 329984 6112
rect 349068 6060 349120 6112
rect 378876 6060 378928 6112
rect 390468 6060 390520 6112
rect 538404 6060 538456 6112
rect 264244 5992 264296 6044
rect 292580 5992 292632 6044
rect 300768 5992 300820 6044
rect 328460 5992 328512 6044
rect 348976 5992 349028 6044
rect 375288 5992 375340 6044
rect 389088 5992 389140 6044
rect 534908 5992 534960 6044
rect 265348 5924 265400 5976
rect 286324 5924 286376 5976
rect 304356 5924 304408 5976
rect 329840 5924 329892 5976
rect 347688 5924 347740 5976
rect 371700 5924 371752 5976
rect 388996 5924 389048 5976
rect 531320 5924 531372 5976
rect 311440 5856 311492 5908
rect 331312 5856 331364 5908
rect 344836 5856 344888 5908
rect 315028 5788 315080 5840
rect 332692 5788 332744 5840
rect 347596 5788 347648 5840
rect 368204 5856 368256 5908
rect 387708 5856 387760 5908
rect 527824 5856 527876 5908
rect 364616 5788 364668 5840
rect 386236 5788 386288 5840
rect 524236 5788 524288 5840
rect 318524 5720 318576 5772
rect 332600 5720 332652 5772
rect 344928 5720 344980 5772
rect 322112 5652 322164 5704
rect 333980 5652 334032 5704
rect 342076 5652 342128 5704
rect 346952 5652 347004 5704
rect 361120 5720 361172 5772
rect 386328 5720 386380 5772
rect 520740 5720 520792 5772
rect 357532 5652 357584 5704
rect 384948 5652 385000 5704
rect 517152 5652 517204 5704
rect 329196 5584 329248 5636
rect 335360 5584 335412 5636
rect 332692 5516 332744 5568
rect 336740 5584 336792 5636
rect 346308 5584 346360 5636
rect 389824 5584 389876 5636
rect 391848 5584 391900 5636
rect 513564 5584 513616 5636
rect 336280 5516 336332 5568
rect 338120 5516 338172 5568
rect 339408 5516 339460 5568
rect 339868 5516 339920 5568
rect 340788 5516 340840 5568
rect 343364 5516 343416 5568
rect 354496 5516 354548 5568
rect 541992 5516 542044 5568
rect 200028 5448 200080 5500
rect 246396 5448 246448 5500
rect 274456 5448 274508 5500
rect 540796 5448 540848 5500
rect 201316 5380 201368 5432
rect 249984 5380 250036 5432
rect 275928 5380 275980 5432
rect 544384 5380 544436 5432
rect 201408 5312 201460 5364
rect 253480 5312 253532 5364
rect 277308 5312 277360 5364
rect 547880 5312 547932 5364
rect 202788 5244 202840 5296
rect 257068 5244 257120 5296
rect 277216 5244 277268 5296
rect 551468 5244 551520 5296
rect 202696 5176 202748 5228
rect 260564 5176 260616 5228
rect 278688 5176 278740 5228
rect 554964 5176 555016 5228
rect 204168 5108 204220 5160
rect 264152 5108 264204 5160
rect 279976 5108 280028 5160
rect 558552 5108 558604 5160
rect 205548 5040 205600 5092
rect 267740 5040 267792 5092
rect 280068 5040 280120 5092
rect 562048 5040 562100 5092
rect 205456 4972 205508 5024
rect 271236 4972 271288 5024
rect 281448 4972 281500 5024
rect 565636 4972 565688 5024
rect 206928 4904 206980 4956
rect 274824 4904 274876 4956
rect 282828 4904 282880 4956
rect 569132 4904 569184 4956
rect 208216 4836 208268 4888
rect 278320 4836 278372 4888
rect 282736 4836 282788 4888
rect 572720 4836 572772 4888
rect 208308 4768 208360 4820
rect 281908 4768 281960 4820
rect 284208 4768 284260 4820
rect 576308 4768 576360 4820
rect 198556 4700 198608 4752
rect 242900 4700 242952 4752
rect 274548 4700 274600 4752
rect 537208 4700 537260 4752
rect 198648 4632 198700 4684
rect 239312 4632 239364 4684
rect 273076 4632 273128 4684
rect 533712 4632 533764 4684
rect 197268 4564 197320 4616
rect 235816 4564 235868 4616
rect 273168 4564 273220 4616
rect 530124 4564 530176 4616
rect 195796 4496 195848 4548
rect 232228 4496 232280 4548
rect 271788 4496 271840 4548
rect 526628 4496 526680 4548
rect 195888 4428 195940 4480
rect 228732 4428 228784 4480
rect 270408 4428 270460 4480
rect 523040 4428 523092 4480
rect 194508 4360 194560 4412
rect 225144 4360 225196 4412
rect 270316 4360 270368 4412
rect 519544 4360 519596 4412
rect 193128 4292 193180 4344
rect 221556 4292 221608 4344
rect 269028 4292 269080 4344
rect 515956 4292 516008 4344
rect 193036 4224 193088 4276
rect 218060 4224 218112 4276
rect 267648 4224 267700 4276
rect 512460 4224 512512 4276
rect 400864 4156 400916 4208
rect 402520 4156 402572 4208
rect 456800 4156 456852 4208
rect 340972 4088 341024 4140
rect 377404 4088 377456 4140
rect 394240 4088 394292 4140
rect 467840 4088 467892 4140
rect 507768 4088 507820 4140
rect 543188 4088 543240 4140
rect 319720 4020 319772 4072
rect 356704 4020 356756 4072
rect 390652 4020 390704 4072
rect 138848 3952 138900 4004
rect 142804 3952 142856 4004
rect 196624 3952 196676 4004
rect 203892 3952 203944 4004
rect 309048 3952 309100 4004
rect 340144 3952 340196 4004
rect 344560 3952 344612 4004
rect 382924 3952 382976 4004
rect 387156 3952 387208 4004
rect 466460 4020 466512 4072
rect 489184 4020 489236 4072
rect 491116 4020 491168 4072
rect 509056 4020 509108 4072
rect 546684 4020 546736 4072
rect 465172 3952 465224 4004
rect 497464 3952 497516 4004
rect 500592 3952 500644 4004
rect 509148 3952 509200 4004
rect 550272 3952 550324 4004
rect 169024 3884 169076 3936
rect 187608 3884 187660 3936
rect 196808 3884 196860 3936
rect 248788 3884 248840 3936
rect 267004 3884 267056 3936
rect 277216 3884 277268 3936
rect 294604 3884 294656 3936
rect 301964 3884 302016 3936
rect 318064 3884 318116 3936
rect 326804 3884 326856 3936
rect 363604 3884 363656 3936
rect 383568 3884 383620 3936
rect 465264 3884 465316 3936
rect 511908 3884 511960 3936
rect 553768 3884 553820 3936
rect 154212 3816 154264 3868
rect 166264 3816 166316 3868
rect 168380 3816 168432 3868
rect 178224 3816 178276 3868
rect 190276 3816 190328 3868
rect 207388 3816 207440 3868
rect 145932 3748 145984 3800
rect 162124 3748 162176 3800
rect 166080 3748 166132 3800
rect 177304 3748 177356 3800
rect 190368 3748 190420 3800
rect 210976 3748 211028 3800
rect 252376 3748 252428 3800
rect 271144 3816 271196 3868
rect 294880 3816 294932 3868
rect 323584 3816 323636 3868
rect 337476 3816 337528 3868
rect 376024 3816 376076 3868
rect 379980 3816 380032 3868
rect 266544 3748 266596 3800
rect 295984 3748 296036 3800
rect 298468 3748 298520 3800
rect 320824 3748 320876 3800
rect 323308 3748 323360 3800
rect 360844 3748 360896 3800
rect 376484 3748 376536 3800
rect 463700 3816 463752 3868
rect 511816 3816 511868 3868
rect 557356 3816 557408 3868
rect 160100 3680 160152 3732
rect 188344 3680 188396 3732
rect 191748 3680 191800 3732
rect 214472 3680 214524 3732
rect 238116 3680 238168 3732
rect 249064 3680 249116 3732
rect 255872 3680 255924 3732
rect 280804 3680 280856 3732
rect 287796 3680 287848 3732
rect 322204 3680 322256 3732
rect 330392 3680 330444 3732
rect 371884 3680 371936 3732
rect 372896 3680 372948 3732
rect 462412 3748 462464 3800
rect 462596 3748 462648 3800
rect 469220 3748 469272 3800
rect 498108 3748 498160 3800
rect 504180 3748 504232 3800
rect 513288 3748 513340 3800
rect 153016 3612 153068 3664
rect 173072 3612 173124 3664
rect 180248 3612 180300 3664
rect 184204 3612 184256 3664
rect 137652 3544 137704 3596
rect 164884 3544 164936 3596
rect 165528 3544 165580 3596
rect 167184 3544 167236 3596
rect 168288 3544 168340 3596
rect 173164 3544 173216 3596
rect 173808 3544 173860 3596
rect 179052 3544 179104 3596
rect 180064 3544 180116 3596
rect 181444 3544 181496 3596
rect 182088 3544 182140 3596
rect 183744 3544 183796 3596
rect 184848 3544 184900 3596
rect 186136 3544 186188 3596
rect 187332 3612 187384 3664
rect 214564 3612 214616 3664
rect 220452 3612 220504 3664
rect 238024 3612 238076 3664
rect 224224 3544 224276 3596
rect 231032 3544 231084 3596
rect 231676 3544 231728 3596
rect 234620 3544 234672 3596
rect 260104 3612 260156 3664
rect 262956 3612 263008 3664
rect 298836 3612 298888 3664
rect 316224 3612 316276 3664
rect 358084 3612 358136 3664
rect 369400 3612 369452 3664
rect 472072 3680 472124 3732
rect 483756 3680 483808 3732
rect 503536 3680 503588 3732
rect 560852 3748 560904 3800
rect 564440 3680 564492 3732
rect 258264 3544 258316 3596
rect 259276 3544 259328 3596
rect 259460 3544 259512 3596
rect 260656 3544 260708 3596
rect 261760 3544 261812 3596
rect 262864 3544 262916 3596
rect 273628 3544 273680 3596
rect 274364 3544 274416 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 278044 3544 278096 3596
rect 280712 3544 280764 3596
rect 318156 3544 318208 3596
rect 333888 3544 333940 3596
rect 334716 3544 334768 3596
rect 340880 3544 340932 3596
rect 342168 3544 342220 3596
rect 351644 3544 351696 3596
rect 454500 3544 454552 3596
rect 455328 3544 455380 3596
rect 458088 3612 458140 3664
rect 484584 3612 484636 3664
rect 498016 3612 498068 3664
rect 507676 3612 507728 3664
rect 514668 3612 514720 3664
rect 568028 3612 568080 3664
rect 462504 3544 462556 3596
rect 467104 3544 467156 3596
rect 510068 3544 510120 3596
rect 510528 3544 510580 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 135260 3476 135312 3528
rect 137284 3476 137336 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 143540 3476 143592 3528
rect 144644 3476 144696 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 150624 3476 150676 3528
rect 151728 3476 151780 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 155408 3476 155460 3528
rect 155868 3476 155920 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 131764 3408 131816 3460
rect 132408 3408 132460 3460
rect 156604 3340 156656 3392
rect 407396 3476 407448 3528
rect 411904 3476 411956 3528
rect 149520 3272 149572 3324
rect 405740 3408 405792 3460
rect 408408 3408 408460 3460
rect 461584 3408 461636 3460
rect 462228 3408 462280 3460
rect 465172 3408 465224 3460
rect 466368 3408 466420 3460
rect 468668 3408 468720 3460
rect 469128 3408 469180 3460
rect 472256 3476 472308 3528
rect 473268 3476 473320 3528
rect 479340 3476 479392 3528
rect 480168 3476 480220 3528
rect 486424 3476 486476 3528
rect 487068 3476 487120 3528
rect 473544 3408 473596 3460
rect 486516 3408 486568 3460
rect 492312 3408 492364 3460
rect 163688 3340 163740 3392
rect 164148 3340 164200 3392
rect 184940 3340 184992 3392
rect 186228 3340 186280 3392
rect 188528 3340 188580 3392
rect 188988 3340 189040 3392
rect 191104 3340 191156 3392
rect 193220 3340 193272 3392
rect 199108 3340 199160 3392
rect 199936 3340 199988 3392
rect 206192 3340 206244 3392
rect 206836 3340 206888 3392
rect 209780 3340 209832 3392
rect 211068 3340 211120 3392
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 216864 3340 216916 3392
rect 217968 3340 218020 3392
rect 241704 3340 241756 3392
rect 242716 3340 242768 3392
rect 245200 3340 245252 3392
rect 246304 3340 246356 3392
rect 254676 3340 254728 3392
rect 255964 3340 256016 3392
rect 270040 3340 270092 3392
rect 305552 3340 305604 3392
rect 306288 3340 306340 3392
rect 312636 3340 312688 3392
rect 342904 3340 342956 3392
rect 348056 3340 348108 3392
rect 378784 3340 378836 3392
rect 397736 3340 397788 3392
rect 460940 3340 460992 3392
rect 467932 3340 467984 3392
rect 489920 3340 489972 3392
rect 491208 3340 491260 3392
rect 493508 3476 493560 3528
rect 493968 3476 494020 3528
rect 504364 3476 504416 3528
rect 505376 3476 505428 3528
rect 507124 3476 507176 3528
rect 508872 3476 508924 3528
rect 514576 3476 514628 3528
rect 571524 3544 571576 3596
rect 516048 3476 516100 3528
rect 575112 3476 575164 3528
rect 493324 3408 493376 3460
rect 494704 3408 494756 3460
rect 500776 3408 500828 3460
rect 514760 3408 514812 3460
rect 517428 3408 517480 3460
rect 578608 3408 578660 3460
rect 499396 3340 499448 3392
rect 499488 3340 499540 3392
rect 511264 3340 511316 3392
rect 162492 3272 162544 3324
rect 170404 3272 170456 3324
rect 192024 3272 192076 3324
rect 192944 3272 192996 3324
rect 223948 3272 224000 3324
rect 228456 3272 228508 3324
rect 401324 3272 401376 3324
rect 470692 3272 470744 3324
rect 495348 3272 495400 3324
rect 497096 3272 497148 3324
rect 506388 3272 506440 3324
rect 283104 3204 283156 3256
rect 284116 3204 284168 3256
rect 404820 3204 404872 3256
rect 470784 3204 470836 3256
rect 506296 3204 506348 3256
rect 539600 3340 539652 3392
rect 536104 3272 536156 3324
rect 141240 3136 141292 3188
rect 142068 3136 142120 3188
rect 175464 3136 175516 3188
rect 178684 3136 178736 3188
rect 291384 3136 291436 3188
rect 298744 3136 298796 3188
rect 422576 3136 422628 3188
rect 423588 3136 423640 3188
rect 186964 3068 187016 3120
rect 189724 3068 189776 3120
rect 418988 3068 419040 3120
rect 474832 3136 474884 3188
rect 505008 3136 505060 3188
rect 532516 3204 532568 3256
rect 529020 3136 529072 3188
rect 174268 3000 174320 3052
rect 175188 3000 175240 3052
rect 284300 3000 284352 3052
rect 285588 3000 285640 3052
rect 415492 3000 415544 3052
rect 416688 3000 416740 3052
rect 426164 3000 426216 3052
rect 476304 3068 476356 3120
rect 503628 3068 503680 3120
rect 525432 3068 525484 3120
rect 429660 3000 429712 3052
rect 477500 3000 477552 3052
rect 490564 3000 490616 3052
rect 498200 3000 498252 3052
rect 502248 3000 502300 3052
rect 521844 3000 521896 3052
rect 171968 2932 172020 2984
rect 179420 2932 179472 2984
rect 440332 2932 440384 2984
rect 441528 2932 441580 2984
rect 447416 2932 447468 2984
rect 448428 2932 448480 2984
rect 436744 2864 436796 2916
rect 478972 2932 479024 2984
rect 500868 2932 500920 2984
rect 518348 2932 518400 2984
rect 443828 2796 443880 2848
rect 481824 2864 481876 2916
rect 450912 2796 450964 2848
rect 483020 2796 483072 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 641714 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3424 641708 3476 641714
rect 3424 641650 3476 641656
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3436 597514 3464 632023
rect 3528 630630 3556 671191
rect 3606 658200 3662 658209
rect 3606 658135 3662 658144
rect 3516 630624 3568 630630
rect 3516 630566 3568 630572
rect 3620 619614 3648 658135
rect 8220 654838 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 702434 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72988 702406 73108 702434
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 654906 24808 699654
rect 41340 654974 41368 700334
rect 41328 654968 41380 654974
rect 41328 654910 41380 654916
rect 24768 654900 24820 654906
rect 24768 654842 24820 654848
rect 73080 654838 73108 702406
rect 89640 654906 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 700398 105492 703520
rect 137848 702434 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137848 702406 137968 702434
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 106200 654974 106228 700334
rect 97540 654968 97592 654974
rect 97540 654910 97592 654916
rect 106188 654968 106240 654974
rect 106188 654910 106240 654916
rect 84752 654900 84804 654906
rect 84752 654842 84804 654848
rect 89628 654900 89680 654906
rect 89628 654842 89680 654848
rect 8208 654832 8260 654838
rect 8208 654774 8260 654780
rect 72976 654832 73028 654838
rect 72976 654774 73028 654780
rect 73068 654832 73120 654838
rect 73068 654774 73120 654780
rect 72988 652202 73016 654774
rect 84764 652202 84792 654842
rect 97552 652202 97580 654910
rect 135996 654900 136048 654906
rect 135996 654842 136048 654848
rect 123116 654832 123168 654838
rect 123116 654774 123168 654780
rect 123128 652202 123156 654774
rect 136008 652202 136036 654842
rect 137940 654838 137968 702406
rect 148784 654968 148836 654974
rect 148784 654910 148836 654916
rect 137928 654832 137980 654838
rect 137928 654774 137980 654780
rect 148796 652202 148824 654910
rect 154500 654906 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 284036 703582 284248 703610
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 171060 654974 171088 700198
rect 171048 654968 171100 654974
rect 171048 654910 171100 654916
rect 199936 654968 199988 654974
rect 199936 654910 199988 654916
rect 154488 654900 154540 654906
rect 154488 654842 154540 654848
rect 187148 654900 187200 654906
rect 187148 654842 187200 654848
rect 174360 654832 174412 654838
rect 174360 654774 174412 654780
rect 174372 652202 174400 654774
rect 187160 652202 187188 654842
rect 199948 652202 199976 654910
rect 202800 654838 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 219360 654906 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 219348 654900 219400 654906
rect 219348 654842 219400 654848
rect 235920 654838 235948 700334
rect 238300 654900 238352 654906
rect 238300 654842 238352 654848
rect 202788 654832 202840 654838
rect 202788 654774 202840 654780
rect 225512 654832 225564 654838
rect 225512 654774 225564 654780
rect 235908 654832 235960 654838
rect 235908 654774 235960 654780
rect 225524 652202 225552 654774
rect 238312 652202 238340 654842
rect 267660 654838 267688 703520
rect 283852 703474 283880 703520
rect 284036 703474 284064 703582
rect 283852 703446 284064 703474
rect 251180 654832 251232 654838
rect 251180 654774 251232 654780
rect 267648 654832 267700 654838
rect 267648 654774 267700 654780
rect 276756 654832 276808 654838
rect 276756 654774 276808 654780
rect 251192 652202 251220 654774
rect 276768 652202 276796 654774
rect 284220 654430 284248 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 699718 300164 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 364996 700330 365024 703520
rect 393228 700392 393280 700398
rect 393228 700334 393280 700340
rect 340788 700324 340840 700330
rect 340788 700266 340840 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 354588 700324 354640 700330
rect 354588 700266 354640 700272
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 379428 700324 379480 700330
rect 379428 700266 379480 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 328368 699712 328420 699718
rect 328368 699654 328420 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 300780 655518 300808 699654
rect 300768 655512 300820 655518
rect 300768 655454 300820 655460
rect 302332 655512 302384 655518
rect 302332 655454 302384 655460
rect 284208 654424 284260 654430
rect 284208 654366 284260 654372
rect 289544 654424 289596 654430
rect 289544 654366 289596 654372
rect 289556 652202 289584 654366
rect 302344 652202 302372 655454
rect 72988 652174 73072 652202
rect 84764 652174 84848 652202
rect 97552 652174 97636 652202
rect 123128 652174 123212 652202
rect 136008 652174 136092 652202
rect 148796 652174 148880 652202
rect 174372 652174 174456 652202
rect 187160 652174 187244 652202
rect 199948 652174 200032 652202
rect 225524 652174 225608 652202
rect 238312 652174 238396 652202
rect 251192 652174 251276 652202
rect 276768 652174 276852 652202
rect 289556 652174 289640 652202
rect 302344 652174 302428 652202
rect 73044 651984 73072 652174
rect 84820 651984 84848 652174
rect 97608 651984 97636 652174
rect 123184 651984 123212 652174
rect 136064 651984 136092 652174
rect 148852 651984 148880 652174
rect 174428 651984 174456 652174
rect 187216 651984 187244 652174
rect 200004 651984 200032 652174
rect 225580 651984 225608 652174
rect 238368 651984 238396 652174
rect 251248 651984 251276 652174
rect 276824 651984 276852 652174
rect 289612 651984 289640 652174
rect 302400 651984 302428 652174
rect 328380 652066 328408 699654
rect 340800 652202 340828 700266
rect 354600 655518 354628 700266
rect 353576 655512 353628 655518
rect 353576 655454 353628 655460
rect 354588 655512 354640 655518
rect 354588 655454 354640 655460
rect 353588 652202 353616 655454
rect 327976 652038 328408 652066
rect 340764 652174 340828 652202
rect 353552 652174 353616 652202
rect 327976 651984 328004 652038
rect 340764 651984 340792 652174
rect 353552 651984 353580 652174
rect 379440 652066 379468 700266
rect 393240 654634 393268 700334
rect 397472 700330 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429856 700330 429884 703520
rect 462332 700466 462360 703520
rect 430488 700460 430540 700466
rect 430488 700402 430540 700408
rect 462320 700460 462372 700466
rect 462320 700402 462372 700408
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 405648 700324 405700 700330
rect 405648 700266 405700 700272
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 405660 654838 405688 700266
rect 404820 654832 404872 654838
rect 404820 654774 404872 654780
rect 405648 654832 405700 654838
rect 405648 654774 405700 654780
rect 392032 654628 392084 654634
rect 392032 654570 392084 654576
rect 393228 654628 393280 654634
rect 393228 654570 393280 654576
rect 392044 652202 392072 654570
rect 404832 652202 404860 654774
rect 379220 652038 379468 652066
rect 392008 652174 392072 652202
rect 404796 652174 404860 652202
rect 379220 651984 379248 652038
rect 392008 651984 392036 652174
rect 404796 651984 404824 652174
rect 430500 652066 430528 700402
rect 478524 700398 478552 703520
rect 482928 700460 482980 700466
rect 482928 700402 482980 700408
rect 444288 700392 444340 700398
rect 444288 700334 444340 700340
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 444300 655518 444328 700334
rect 456708 700324 456760 700330
rect 456708 700266 456760 700272
rect 456720 655518 456748 700266
rect 482940 655518 482968 700402
rect 494808 700330 494836 703520
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 495348 700392 495400 700398
rect 495348 700334 495400 700340
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 443184 655512 443236 655518
rect 443184 655454 443236 655460
rect 444288 655512 444340 655518
rect 444288 655454 444340 655460
rect 455972 655512 456024 655518
rect 455972 655454 456024 655460
rect 456708 655512 456760 655518
rect 456708 655454 456760 655460
rect 481640 655512 481692 655518
rect 481640 655454 481692 655460
rect 482928 655512 482980 655518
rect 482928 655454 482980 655460
rect 443196 652202 443224 655454
rect 455984 652202 456012 655454
rect 481652 652202 481680 655454
rect 495360 655042 495388 700334
rect 559668 700330 559696 703520
rect 507768 700324 507820 700330
rect 507768 700266 507820 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 494428 655036 494480 655042
rect 494428 654978 494480 654984
rect 495348 655036 495400 655042
rect 495348 654978 495400 654984
rect 494440 652202 494468 654978
rect 507780 654430 507808 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 522304 696992 522356 696998
rect 522304 696934 522356 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 507216 654424 507268 654430
rect 507216 654366 507268 654372
rect 507768 654424 507820 654430
rect 507768 654366 507820 654372
rect 507228 652202 507256 654366
rect 430372 652038 430528 652066
rect 443160 652174 443224 652202
rect 455948 652174 456012 652202
rect 481616 652174 481680 652202
rect 494404 652174 494468 652202
rect 507192 652174 507256 652202
rect 430372 651984 430400 652038
rect 443160 651984 443188 652174
rect 455948 651984 455976 652174
rect 481616 651984 481644 652174
rect 494404 651984 494432 652174
rect 507192 651984 507220 652174
rect 522316 650865 522344 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 522396 683188 522448 683194
rect 522396 683130 522448 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 522302 650856 522358 650865
rect 522302 650791 522358 650800
rect 522304 643136 522356 643142
rect 522304 643078 522356 643084
rect 69020 641708 69072 641714
rect 69020 641650 69072 641656
rect 69032 640937 69060 641650
rect 69018 640928 69074 640937
rect 69018 640863 69074 640872
rect 69020 630624 69072 630630
rect 69020 630566 69072 630572
rect 69032 629785 69060 630566
rect 69018 629776 69074 629785
rect 69018 629711 69074 629720
rect 3608 619608 3660 619614
rect 3608 619550 3660 619556
rect 69020 619608 69072 619614
rect 69020 619550 69072 619556
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 597508 3476 597514
rect 3424 597450 3476 597456
rect 3528 585138 3556 619103
rect 69032 618633 69060 619550
rect 69018 618624 69074 618633
rect 69018 618559 69074 618568
rect 522316 606529 522344 643078
rect 522408 640529 522436 683130
rect 522488 670744 522540 670750
rect 580172 670744 580224 670750
rect 522488 670686 522540 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 522394 640520 522450 640529
rect 522394 640455 522450 640464
rect 522396 630692 522448 630698
rect 522396 630634 522448 630640
rect 522302 606520 522358 606529
rect 522302 606455 522358 606464
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3516 585132 3568 585138
rect 3516 585074 3568 585080
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 552022 3464 579935
rect 3620 574054 3648 606047
rect 69020 597508 69072 597514
rect 69020 597450 69072 597456
rect 69032 596329 69060 597450
rect 69018 596320 69074 596329
rect 69018 596255 69074 596264
rect 522408 595105 522436 630634
rect 522500 629241 522528 670686
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 522486 629232 522542 629241
rect 522486 629167 522542 629176
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 522488 616888 522540 616894
rect 522488 616830 522540 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 522394 595096 522450 595105
rect 522394 595031 522450 595040
rect 522304 590708 522356 590714
rect 522304 590650 522356 590656
rect 69020 585132 69072 585138
rect 69020 585074 69072 585080
rect 69032 585041 69060 585074
rect 69018 585032 69074 585041
rect 69018 584967 69074 584976
rect 3608 574048 3660 574054
rect 3608 573990 3660 573996
rect 69020 574048 69072 574054
rect 69020 573990 69072 573996
rect 69032 573889 69060 573990
rect 69018 573880 69074 573889
rect 69018 573815 69074 573824
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 552016 3476 552022
rect 3424 551958 3476 551964
rect 3528 540938 3556 566879
rect 522316 560833 522344 590650
rect 522500 583681 522528 616830
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 522486 583672 522542 583681
rect 522486 583607 522542 583616
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 522396 576904 522448 576910
rect 522396 576846 522448 576852
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 522302 560824 522358 560833
rect 522302 560759 522358 560768
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3516 540932 3568 540938
rect 3516 540874 3568 540880
rect 3620 529922 3648 553823
rect 69020 552016 69072 552022
rect 69020 551958 69072 551964
rect 69032 551585 69060 551958
rect 69018 551576 69074 551585
rect 69018 551511 69074 551520
rect 522408 549545 522436 576846
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 522488 563100 522540 563106
rect 522488 563042 522540 563048
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 522394 549536 522450 549545
rect 522394 549471 522450 549480
rect 69020 540932 69072 540938
rect 69020 540874 69072 540880
rect 69032 540433 69060 540874
rect 69018 540424 69074 540433
rect 69018 540359 69074 540368
rect 522500 538121 522528 563042
rect 522486 538112 522542 538121
rect 522486 538047 522542 538056
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 522304 536852 522356 536858
rect 522304 536794 522356 536800
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 3608 529916 3660 529922
rect 3608 529858 3660 529864
rect 69020 529916 69072 529922
rect 69020 529858 69072 529864
rect 69032 529281 69060 529858
rect 69018 529272 69074 529281
rect 69018 529207 69074 529216
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 507822 3464 527847
rect 522316 515409 522344 536794
rect 580170 524512 580226 524521
rect 522396 524476 522448 524482
rect 580170 524447 580172 524456
rect 522396 524418 522448 524424
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 522302 515400 522358 515409
rect 522302 515335 522358 515344
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 507816 3476 507822
rect 3424 507758 3476 507764
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3436 485790 3464 501735
rect 3528 496806 3556 514791
rect 522304 510672 522356 510678
rect 522304 510614 522356 510620
rect 69020 507816 69072 507822
rect 69020 507758 69072 507764
rect 69032 506977 69060 507758
rect 69018 506968 69074 506977
rect 69018 506903 69074 506912
rect 3516 496800 3568 496806
rect 3516 496742 3568 496748
rect 69020 496800 69072 496806
rect 69020 496742 69072 496748
rect 69032 495689 69060 496742
rect 69018 495680 69074 495689
rect 69018 495615 69074 495624
rect 522316 492561 522344 510614
rect 522408 503985 522436 524418
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 522394 503976 522450 503985
rect 522394 503911 522450 503920
rect 522302 492552 522358 492561
rect 522302 492487 522358 492496
rect 3424 485784 3476 485790
rect 3424 485726 3476 485732
rect 69020 485784 69072 485790
rect 69020 485726 69072 485732
rect 69032 484537 69060 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 69018 484528 69074 484537
rect 69018 484463 69074 484472
rect 580184 484430 580212 484599
rect 522304 484424 522356 484430
rect 522304 484366 522356 484372
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 462330 3464 475623
rect 522316 469849 522344 484366
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 522396 470620 522448 470626
rect 522396 470562 522448 470568
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 522302 469840 522358 469849
rect 522302 469775 522358 469784
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3424 462324 3476 462330
rect 3424 462266 3476 462272
rect 3528 451246 3556 462567
rect 69020 462324 69072 462330
rect 69020 462266 69072 462272
rect 69032 462233 69060 462266
rect 69018 462224 69074 462233
rect 69018 462159 69074 462168
rect 522408 458425 522436 470562
rect 522394 458416 522450 458425
rect 522394 458351 522450 458360
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 522304 456816 522356 456822
rect 522304 456758 522356 456764
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 3516 451240 3568 451246
rect 3516 451182 3568 451188
rect 69020 451240 69072 451246
rect 69020 451182 69072 451188
rect 69032 451081 69060 451182
rect 69018 451072 69074 451081
rect 69018 451007 69074 451016
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3436 440230 3464 449511
rect 522316 447001 522344 456758
rect 522302 446992 522358 447001
rect 522302 446927 522358 446936
rect 3424 440224 3476 440230
rect 3424 440166 3476 440172
rect 69020 440224 69072 440230
rect 69020 440166 69072 440172
rect 69032 439929 69060 440166
rect 69018 439920 69074 439929
rect 69018 439855 69074 439864
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 522948 430636 523000 430642
rect 522948 430578 523000 430584
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 522960 424289 522988 430578
rect 522946 424280 523002 424289
rect 522946 424215 523002 424224
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 418130 3372 423535
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 522948 418192 523000 418198
rect 522948 418134 523000 418140
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 3332 418124 3384 418130
rect 3332 418066 3384 418072
rect 69020 418124 69072 418130
rect 69020 418066 69072 418072
rect 69032 417489 69060 418066
rect 69018 417480 69074 417489
rect 69018 417415 69074 417424
rect 522960 412865 522988 418134
rect 522946 412856 523002 412865
rect 522946 412791 523002 412800
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 407114 3464 410479
rect 3424 407108 3476 407114
rect 3424 407050 3476 407056
rect 69020 407108 69072 407114
rect 69020 407050 69072 407056
rect 69032 406473 69060 407050
rect 69018 406464 69074 406473
rect 69018 406399 69074 406408
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 522028 404388 522080 404394
rect 522028 404330 522080 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 522040 401577 522068 404330
rect 522026 401568 522082 401577
rect 522026 401503 522082 401512
rect 2870 397488 2926 397497
rect 2870 397423 2926 397432
rect 2884 396030 2912 397423
rect 2872 396024 2924 396030
rect 2872 395966 2924 395972
rect 69020 396024 69072 396030
rect 69020 395966 69072 395972
rect 69032 395185 69060 395966
rect 69018 395176 69074 395185
rect 69018 395111 69074 395120
rect 522948 378820 523000 378826
rect 522948 378762 523000 378768
rect 580172 378820 580224 378826
rect 580172 378762 580224 378768
rect 522960 378729 522988 378762
rect 522946 378720 523002 378729
rect 522946 378655 523002 378664
rect 580184 378457 580212 378762
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 69018 372872 69074 372881
rect 69018 372807 69074 372816
rect 69032 372638 69060 372807
rect 3424 372632 3476 372638
rect 3424 372574 3476 372580
rect 69020 372632 69072 372638
rect 69020 372574 69072 372580
rect 3436 371385 3464 372574
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 522946 367296 523002 367305
rect 522946 367231 523002 367240
rect 522960 365702 522988 367231
rect 522948 365696 523000 365702
rect 522948 365638 523000 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 69018 361720 69074 361729
rect 69018 361655 69074 361664
rect 69032 361622 69060 361655
rect 3424 361616 3476 361622
rect 3424 361558 3476 361564
rect 69020 361616 69072 361622
rect 69020 361558 69072 361564
rect 3436 358465 3464 361558
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 522946 356008 523002 356017
rect 522946 355943 523002 355952
rect 522960 353258 522988 355943
rect 522948 353252 523000 353258
rect 522948 353194 523000 353200
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 69018 350432 69074 350441
rect 69018 350367 69074 350376
rect 69032 349178 69060 350367
rect 2872 349172 2924 349178
rect 2872 349114 2924 349120
rect 69020 349172 69072 349178
rect 69020 349114 69072 349120
rect 2884 345409 2912 349114
rect 2870 345400 2926 345409
rect 2870 345335 2926 345344
rect 522302 333160 522358 333169
rect 522302 333095 522358 333104
rect 69018 328128 69074 328137
rect 69018 328063 69074 328072
rect 69032 327146 69060 328063
rect 2872 327140 2924 327146
rect 2872 327082 2924 327088
rect 69020 327140 69072 327146
rect 69020 327082 69072 327088
rect 2884 319297 2912 327082
rect 522316 325650 522344 333095
rect 522304 325644 522356 325650
rect 522304 325586 522356 325592
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 522302 321872 522358 321881
rect 522302 321807 522358 321816
rect 2870 319288 2926 319297
rect 2870 319223 2926 319232
rect 69018 316976 69074 316985
rect 69018 316911 69074 316920
rect 69032 316062 69060 316911
rect 3516 316056 3568 316062
rect 3516 315998 3568 316004
rect 69020 316056 69072 316062
rect 69020 315998 69072 316004
rect 3528 306241 3556 315998
rect 522316 313274 522344 321807
rect 522304 313268 522356 313274
rect 522304 313210 522356 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 522302 310312 522358 310321
rect 522302 310247 522358 310256
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 69018 305824 69074 305833
rect 69018 305759 69074 305768
rect 69032 305046 69060 305759
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 69020 305040 69072 305046
rect 69020 304982 69072 304988
rect 3436 293185 3464 304982
rect 522316 299470 522344 310247
rect 522304 299464 522356 299470
rect 522304 299406 522356 299412
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 522394 287736 522450 287745
rect 522394 287671 522450 287680
rect 69018 283384 69074 283393
rect 69018 283319 69074 283328
rect 69032 282946 69060 283319
rect 3424 282940 3476 282946
rect 3424 282882 3476 282888
rect 69020 282940 69072 282946
rect 69020 282882 69072 282888
rect 3436 267209 3464 282882
rect 522302 276176 522358 276185
rect 522302 276111 522358 276120
rect 69018 272368 69074 272377
rect 69018 272303 69074 272312
rect 69032 271930 69060 272303
rect 3516 271924 3568 271930
rect 3516 271866 3568 271872
rect 69020 271924 69072 271930
rect 69020 271866 69072 271872
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3424 260908 3476 260914
rect 3424 260850 3476 260856
rect 3436 241097 3464 260850
rect 3528 254153 3556 271866
rect 69018 261080 69074 261089
rect 69018 261015 69074 261024
rect 69032 260914 69060 261015
rect 69020 260908 69072 260914
rect 69020 260850 69072 260856
rect 522316 259418 522344 276111
rect 522408 273222 522436 287671
rect 522396 273216 522448 273222
rect 522396 273158 522448 273164
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 522394 264888 522450 264897
rect 522394 264823 522450 264832
rect 522304 259412 522356 259418
rect 522304 259354 522356 259360
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 522302 253464 522358 253473
rect 522302 253399 522358 253408
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3516 238808 3568 238814
rect 69020 238808 69072 238814
rect 3516 238750 3568 238756
rect 69018 238776 69020 238785
rect 69072 238776 69074 238785
rect 3424 215348 3476 215354
rect 3424 215290 3476 215296
rect 3436 188873 3464 215290
rect 3528 214985 3556 238750
rect 69018 238711 69074 238720
rect 522316 233238 522344 253399
rect 522408 245614 522436 264823
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 522396 245608 522448 245614
rect 580172 245608 580224 245614
rect 522396 245550 522448 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 522394 242040 522450 242049
rect 522394 241975 522450 241984
rect 522304 233232 522356 233238
rect 522304 233174 522356 233180
rect 522302 230752 522358 230761
rect 522302 230687 522358 230696
rect 69018 227624 69074 227633
rect 69018 227559 69074 227568
rect 69032 226370 69060 227559
rect 3608 226364 3660 226370
rect 3608 226306 3660 226312
rect 69020 226364 69072 226370
rect 69020 226306 69072 226312
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3620 201929 3648 226306
rect 69018 216472 69074 216481
rect 69018 216407 69074 216416
rect 69032 215354 69060 216407
rect 69020 215348 69072 215354
rect 69020 215290 69072 215296
rect 522316 206990 522344 230687
rect 522408 219434 522436 241975
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 522396 219428 522448 219434
rect 522396 219370 522448 219376
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 522486 219328 522542 219337
rect 522486 219263 522542 219272
rect 522394 207904 522450 207913
rect 522394 207839 522450 207848
rect 522304 206984 522356 206990
rect 522304 206926 522356 206932
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 522302 196480 522358 196489
rect 522302 196415 522358 196424
rect 69018 194168 69074 194177
rect 69018 194103 69074 194112
rect 69032 193254 69060 194103
rect 3608 193248 3660 193254
rect 3608 193190 3660 193196
rect 69020 193248 69072 193254
rect 69020 193190 69072 193196
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3516 182232 3568 182238
rect 3516 182174 3568 182180
rect 3424 171148 3476 171154
rect 3424 171090 3476 171096
rect 3436 136785 3464 171090
rect 3528 149841 3556 182174
rect 3620 162897 3648 193190
rect 69018 182880 69074 182889
rect 69018 182815 69074 182824
rect 69032 182238 69060 182815
rect 69020 182232 69072 182238
rect 69020 182174 69072 182180
rect 69018 171728 69074 171737
rect 69018 171663 69074 171672
rect 69032 171154 69060 171663
rect 69020 171148 69072 171154
rect 69020 171090 69072 171096
rect 522316 167006 522344 196415
rect 522408 179382 522436 207839
rect 522500 193186 522528 219263
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 522488 193180 522540 193186
rect 522488 193122 522540 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 522486 185192 522542 185201
rect 522486 185127 522542 185136
rect 522396 179376 522448 179382
rect 522396 179318 522448 179324
rect 522394 173904 522450 173913
rect 522394 173839 522450 173848
rect 522304 167000 522356 167006
rect 522304 166942 522356 166948
rect 3606 162888 3662 162897
rect 3606 162823 3662 162832
rect 522302 162344 522358 162353
rect 522302 162279 522358 162288
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 69018 149424 69074 149433
rect 69018 149359 69074 149368
rect 69032 149122 69060 149359
rect 3700 149116 3752 149122
rect 3700 149058 3752 149064
rect 69020 149116 69072 149122
rect 69020 149058 69072 149064
rect 3608 138032 3660 138038
rect 3608 137974 3660 137980
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3516 127016 3568 127022
rect 3516 126958 3568 126964
rect 3424 114572 3476 114578
rect 3424 114514 3476 114520
rect 3436 71641 3464 114514
rect 3528 84697 3556 126958
rect 3620 97617 3648 137974
rect 3712 110673 3740 149058
rect 69018 138272 69074 138281
rect 69018 138207 69074 138216
rect 69032 138038 69060 138207
rect 69020 138032 69072 138038
rect 69020 137974 69072 137980
rect 69018 127120 69074 127129
rect 69018 127055 69074 127064
rect 69032 127022 69060 127055
rect 69020 127016 69072 127022
rect 69020 126958 69072 126964
rect 522316 126954 522344 162279
rect 522408 139398 522436 173839
rect 522500 153202 522528 185127
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 522488 153196 522540 153202
rect 522488 153138 522540 153144
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 522578 151056 522634 151065
rect 522578 150991 522634 151000
rect 522486 139632 522542 139641
rect 522486 139567 522542 139576
rect 522396 139392 522448 139398
rect 522396 139334 522448 139340
rect 522394 128208 522450 128217
rect 522394 128143 522450 128152
rect 522304 126948 522356 126954
rect 522304 126890 522356 126896
rect 522302 116920 522358 116929
rect 522302 116855 522358 116864
rect 69018 115832 69074 115841
rect 69018 115767 69074 115776
rect 69032 114578 69060 115767
rect 69020 114572 69072 114578
rect 69020 114514 69072 114520
rect 3698 110664 3754 110673
rect 3698 110599 3754 110608
rect 69018 104816 69074 104825
rect 69018 104751 69074 104760
rect 69032 103562 69060 104751
rect 3792 103556 3844 103562
rect 3792 103498 3844 103504
rect 69020 103556 69072 103562
rect 69020 103498 69072 103504
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3700 92540 3752 92546
rect 3700 92482 3752 92488
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3608 81456 3660 81462
rect 3608 81398 3660 81404
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3516 70440 3568 70446
rect 3516 70382 3568 70388
rect 3424 60784 3476 60790
rect 3424 60726 3476 60732
rect 2688 57384 2740 57390
rect 2688 57326 2740 57332
rect 1308 57248 1360 57254
rect 1308 57190 1360 57196
rect 1320 3534 1348 57190
rect 2700 3534 2728 57326
rect 3436 6497 3464 60726
rect 3528 19417 3556 70382
rect 3620 32473 3648 81398
rect 3712 45529 3740 92482
rect 3804 58585 3832 103498
rect 69018 93528 69074 93537
rect 69018 93463 69074 93472
rect 69032 92546 69060 93463
rect 69020 92540 69072 92546
rect 69020 92482 69072 92488
rect 69018 82376 69074 82385
rect 69018 82311 69074 82320
rect 69032 81462 69060 82311
rect 69020 81456 69072 81462
rect 69020 81398 69072 81404
rect 522316 73166 522344 116855
rect 522408 86970 522436 128143
rect 522500 100706 522528 139567
rect 522592 113150 522620 150991
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 522580 113144 522632 113150
rect 522580 113086 522632 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 522670 105496 522726 105505
rect 522670 105431 522726 105440
rect 522488 100700 522540 100706
rect 522488 100642 522540 100648
rect 522578 94072 522634 94081
rect 522578 94007 522634 94016
rect 522396 86964 522448 86970
rect 522396 86906 522448 86912
rect 522486 82784 522542 82793
rect 522486 82719 522542 82728
rect 522304 73160 522356 73166
rect 522304 73102 522356 73108
rect 522394 71360 522450 71369
rect 522394 71295 522450 71304
rect 69018 71224 69074 71233
rect 69018 71159 69074 71168
rect 69032 70446 69060 71159
rect 69020 70440 69072 70446
rect 69020 70382 69072 70388
rect 69018 61160 69074 61169
rect 69018 61095 69074 61104
rect 69032 60790 69060 61095
rect 522302 60888 522358 60897
rect 522302 60823 522358 60832
rect 69020 60784 69072 60790
rect 69020 60726 69072 60732
rect 72860 59786 72888 60044
rect 72804 59758 72888 59786
rect 72952 59786 72980 60044
rect 168264 59786 168292 60044
rect 169184 59786 169212 60044
rect 170104 59786 170132 60044
rect 170932 59786 170960 60044
rect 171852 59786 171880 60044
rect 172772 59786 172800 60044
rect 173692 59786 173720 60044
rect 174612 59786 174640 60044
rect 175532 59786 175560 60044
rect 176452 59786 176480 60044
rect 177372 59786 177400 60044
rect 178292 59922 178320 60044
rect 72952 59758 73016 59786
rect 3790 58576 3846 58585
rect 3790 58511 3846 58520
rect 72804 57390 72832 59758
rect 72792 57384 72844 57390
rect 72792 57326 72844 57332
rect 72988 57254 73016 59758
rect 168208 59758 168292 59786
rect 169128 59758 169212 59786
rect 170048 59758 170132 59786
rect 170876 59758 170960 59786
rect 171796 59758 171880 59786
rect 172716 59758 172800 59786
rect 173636 59758 173720 59786
rect 174556 59758 174640 59786
rect 175476 59758 175560 59786
rect 176396 59758 176480 59786
rect 177316 59758 177400 59786
rect 178144 59894 178320 59922
rect 155868 57928 155920 57934
rect 155868 57870 155920 57876
rect 153108 57860 153160 57866
rect 153108 57802 153160 57808
rect 136548 57792 136600 57798
rect 136548 57734 136600 57740
rect 133788 57452 133840 57458
rect 133788 57394 133840 57400
rect 129648 57384 129700 57390
rect 129648 57326 129700 57332
rect 126888 57316 126940 57322
rect 126888 57258 126940 57264
rect 72976 57248 73028 57254
rect 72976 57190 73028 57196
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 126900 3534 126928 57258
rect 128176 10328 128228 10334
rect 128176 10270 128228 10276
rect 126980 7064 127032 7070
rect 126980 7006 127032 7012
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 125888 480 125916 3470
rect 126992 480 127020 7006
rect 128188 480 128216 10270
rect 129660 6914 129688 57326
rect 132408 10396 132460 10402
rect 132408 10338 132460 10344
rect 130568 8968 130620 8974
rect 130568 8910 130620 8916
rect 129384 6886 129688 6914
rect 129384 480 129412 6886
rect 130580 480 130608 8910
rect 132420 3466 132448 10338
rect 133800 3534 133828 57394
rect 134156 9036 134208 9042
rect 134156 8978 134208 8984
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 132408 3460 132460 3466
rect 132408 3402 132460 3408
rect 131776 480 131804 3402
rect 132972 480 133000 3470
rect 134168 480 134196 8978
rect 136560 6914 136588 57734
rect 148968 57724 149020 57730
rect 148968 57666 149020 57672
rect 144828 57656 144880 57662
rect 144828 57598 144880 57604
rect 142068 57588 142120 57594
rect 142068 57530 142120 57536
rect 140688 57520 140740 57526
rect 140688 57462 140740 57468
rect 137284 55888 137336 55894
rect 137284 55830 137336 55836
rect 136468 6886 136588 6914
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 135272 480 135300 3470
rect 136468 480 136496 6886
rect 137296 3534 137324 55830
rect 138848 4004 138900 4010
rect 138848 3946 138900 3952
rect 137652 3596 137704 3602
rect 137652 3538 137704 3544
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 137664 480 137692 3538
rect 138860 480 138888 3946
rect 140700 3534 140728 57462
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 140056 480 140084 3470
rect 142080 3194 142108 57530
rect 144736 57112 144788 57118
rect 144736 57054 144788 57060
rect 143448 54528 143500 54534
rect 143448 54470 143500 54476
rect 142804 28280 142856 28286
rect 142804 28222 142856 28228
rect 142816 4010 142844 28222
rect 142804 4004 142856 4010
rect 142804 3946 142856 3952
rect 143460 3534 143488 54470
rect 144748 16574 144776 57054
rect 144656 16546 144776 16574
rect 144656 3534 144684 16546
rect 144840 6914 144868 57598
rect 147588 56976 147640 56982
rect 147588 56918 147640 56924
rect 144748 6886 144868 6914
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144644 3528 144696 3534
rect 144644 3470 144696 3476
rect 141240 3188 141292 3194
rect 141240 3130 141292 3136
rect 142068 3188 142120 3194
rect 142068 3130 142120 3136
rect 141252 480 141280 3130
rect 142448 480 142476 3470
rect 143552 480 143580 3470
rect 144748 480 144776 6886
rect 145932 3800 145984 3806
rect 145932 3742 145984 3748
rect 145944 480 145972 3742
rect 147600 3534 147628 56918
rect 148980 3534 149008 57666
rect 151728 57044 151780 57050
rect 151728 56986 151780 56992
rect 151740 3534 151768 56986
rect 153016 3664 153068 3670
rect 153016 3606 153068 3612
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149520 3324 149572 3330
rect 149520 3266 149572 3272
rect 149532 480 149560 3266
rect 150636 480 150664 3470
rect 151832 480 151860 3470
rect 153028 480 153056 3606
rect 153120 3534 153148 57802
rect 154212 3868 154264 3874
rect 154212 3810 154264 3816
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154224 480 154252 3810
rect 155880 3534 155908 57870
rect 168208 57322 168236 59758
rect 169128 57390 169156 59758
rect 170048 57458 170076 59758
rect 170876 57798 170904 59758
rect 170864 57792 170916 57798
rect 170864 57734 170916 57740
rect 171796 57526 171824 59758
rect 171784 57520 171836 57526
rect 171784 57462 171836 57468
rect 170036 57452 170088 57458
rect 170036 57394 170088 57400
rect 169116 57384 169168 57390
rect 169116 57326 169168 57332
rect 168196 57316 168248 57322
rect 168196 57258 168248 57264
rect 162124 57248 162176 57254
rect 162124 57190 162176 57196
rect 158628 56908 158680 56914
rect 158628 56850 158680 56856
rect 158640 3534 158668 56850
rect 161388 56840 161440 56846
rect 161388 56782 161440 56788
rect 160008 54596 160060 54602
rect 160008 54538 160060 54544
rect 160020 3534 160048 54538
rect 161400 6914 161428 56782
rect 161308 6886 161428 6914
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 155408 3528 155460 3534
rect 155408 3470 155460 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 155420 480 155448 3470
rect 156604 3392 156656 3398
rect 156604 3334 156656 3340
rect 156616 480 156644 3334
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3674
rect 161308 480 161336 6886
rect 162136 3806 162164 57190
rect 169024 57180 169076 57186
rect 169024 57122 169076 57128
rect 165528 56772 165580 56778
rect 165528 56714 165580 56720
rect 164148 10464 164200 10470
rect 164148 10406 164200 10412
rect 162124 3800 162176 3806
rect 162124 3742 162176 3748
rect 164160 3398 164188 10406
rect 165540 3602 165568 56714
rect 166264 56704 166316 56710
rect 166264 56646 166316 56652
rect 166276 3874 166304 56646
rect 168288 10532 168340 10538
rect 168288 10474 168340 10480
rect 166264 3868 166316 3874
rect 166264 3810 166316 3816
rect 166080 3800 166132 3806
rect 166080 3742 166132 3748
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 165528 3596 165580 3602
rect 165528 3538 165580 3544
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 162492 3324 162544 3330
rect 162492 3266 162544 3272
rect 162504 480 162532 3266
rect 163700 480 163728 3334
rect 164896 480 164924 3538
rect 166092 480 166120 3742
rect 168300 3602 168328 10474
rect 169036 3942 169064 57122
rect 172716 57118 172744 59758
rect 173164 57316 173216 57322
rect 173164 57258 173216 57264
rect 172704 57112 172756 57118
rect 172704 57054 172756 57060
rect 170404 56160 170456 56166
rect 170404 56102 170456 56108
rect 169668 25560 169720 25566
rect 169668 25502 169720 25508
rect 169680 6914 169708 25502
rect 169588 6886 169708 6914
rect 169024 3936 169076 3942
rect 169024 3878 169076 3884
rect 168380 3868 168432 3874
rect 168380 3810 168432 3816
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 168288 3596 168340 3602
rect 168288 3538 168340 3544
rect 167196 480 167224 3538
rect 168392 480 168420 3810
rect 169588 480 169616 6886
rect 170416 3330 170444 56102
rect 170772 10600 170824 10606
rect 170772 10542 170824 10548
rect 170404 3324 170456 3330
rect 170404 3266 170456 3272
rect 170784 480 170812 10542
rect 173176 6914 173204 57258
rect 173636 56982 173664 59758
rect 174556 57050 174584 59758
rect 174544 57044 174596 57050
rect 174544 56986 174596 56992
rect 173624 56976 173676 56982
rect 173624 56918 173676 56924
rect 175476 56710 175504 59758
rect 176396 56914 176424 59758
rect 176384 56908 176436 56914
rect 176384 56850 176436 56856
rect 177316 56846 177344 59758
rect 177304 56840 177356 56846
rect 177304 56782 177356 56788
rect 178144 56778 178172 59894
rect 179120 59786 179148 60044
rect 180040 59786 180068 60044
rect 180960 59786 180988 60044
rect 181880 59786 181908 60044
rect 182800 59786 182828 60044
rect 178236 59758 179148 59786
rect 179432 59758 180068 59786
rect 180904 59758 180988 59786
rect 181824 59758 181908 59786
rect 182192 59758 182828 59786
rect 183720 59786 183748 60044
rect 184640 59786 184668 60044
rect 185560 59786 185588 60044
rect 186388 59786 186416 60044
rect 187308 59786 187336 60044
rect 188228 59786 188256 60044
rect 189148 59786 189176 60044
rect 190068 59786 190096 60044
rect 190988 59786 191016 60044
rect 191908 59786 191936 60044
rect 192828 59786 192856 60044
rect 193656 59786 193684 60044
rect 194576 59786 194604 60044
rect 195496 59786 195524 60044
rect 196416 59786 196444 60044
rect 197336 59786 197364 60044
rect 198256 59786 198284 60044
rect 199176 59786 199204 60044
rect 200096 59786 200124 60044
rect 200924 59786 200952 60044
rect 201844 59786 201872 60044
rect 202764 59786 202792 60044
rect 183720 59758 183784 59786
rect 184640 59758 184704 59786
rect 185560 59758 185624 59786
rect 186388 59758 186452 59786
rect 187308 59758 187372 59786
rect 188228 59758 188292 59786
rect 189148 59758 189212 59786
rect 190068 59758 190408 59786
rect 190988 59758 191052 59786
rect 191908 59758 191972 59786
rect 192828 59758 193168 59786
rect 193656 59758 193720 59786
rect 194576 59758 194640 59786
rect 195496 59758 195836 59786
rect 196416 59758 196480 59786
rect 197336 59758 197400 59786
rect 198256 59758 198596 59786
rect 199176 59758 199240 59786
rect 200096 59758 200160 59786
rect 200924 59758 200988 59786
rect 201844 59758 201908 59786
rect 178132 56772 178184 56778
rect 178132 56714 178184 56720
rect 175464 56704 175516 56710
rect 175464 56646 175516 56652
rect 177304 56228 177356 56234
rect 177304 56170 177356 56176
rect 173808 14884 173860 14890
rect 173808 14826 173860 14832
rect 173084 6886 173204 6914
rect 173084 3670 173112 6886
rect 173072 3664 173124 3670
rect 173072 3606 173124 3612
rect 173820 3602 173848 14826
rect 175188 10668 175240 10674
rect 175188 10610 175240 10616
rect 173164 3596 173216 3602
rect 173164 3538 173216 3544
rect 173808 3596 173860 3602
rect 173808 3538 173860 3544
rect 171968 2984 172020 2990
rect 171968 2926 172020 2932
rect 171980 480 172008 2926
rect 173176 480 173204 3538
rect 175200 3058 175228 10610
rect 176660 6588 176712 6594
rect 176660 6530 176712 6536
rect 175464 3188 175516 3194
rect 175464 3130 175516 3136
rect 174268 3052 174320 3058
rect 174268 2994 174320 3000
rect 175188 3052 175240 3058
rect 175188 2994 175240 3000
rect 174280 480 174308 2994
rect 175476 480 175504 3130
rect 176672 480 176700 6530
rect 177316 3806 177344 56170
rect 177856 10736 177908 10742
rect 177856 10678 177908 10684
rect 177304 3800 177356 3806
rect 177304 3742 177356 3748
rect 177868 480 177896 10678
rect 178236 3874 178264 59758
rect 178684 56704 178736 56710
rect 178684 56646 178736 56652
rect 178224 3868 178276 3874
rect 178224 3810 178276 3816
rect 178696 3194 178724 56646
rect 179052 3596 179104 3602
rect 179052 3538 179104 3544
rect 178684 3188 178736 3194
rect 178684 3130 178736 3136
rect 179064 480 179092 3538
rect 179432 2990 179460 59758
rect 180904 56710 180932 59758
rect 180892 56704 180944 56710
rect 180892 56646 180944 56652
rect 181824 56642 181852 59758
rect 180064 56636 180116 56642
rect 180064 56578 180116 56584
rect 181812 56636 181864 56642
rect 181812 56578 181864 56584
rect 180076 3602 180104 56578
rect 182088 10804 182140 10810
rect 182088 10746 182140 10752
rect 180248 3664 180300 3670
rect 180248 3606 180300 3612
rect 180064 3596 180116 3602
rect 180064 3538 180116 3544
rect 179420 2984 179472 2990
rect 179420 2926 179472 2932
rect 180260 480 180288 3606
rect 182100 3602 182128 10746
rect 181444 3596 181496 3602
rect 181444 3538 181496 3544
rect 182088 3596 182140 3602
rect 182088 3538 182140 3544
rect 181456 480 181484 3538
rect 182192 490 182220 59758
rect 183756 57526 183784 59758
rect 184676 57798 184704 59758
rect 184664 57792 184716 57798
rect 184664 57734 184716 57740
rect 183744 57520 183796 57526
rect 183744 57462 183796 57468
rect 184848 57520 184900 57526
rect 184848 57462 184900 57468
rect 184204 35216 184256 35222
rect 184204 35158 184256 35164
rect 184216 3670 184244 35158
rect 184204 3664 184256 3670
rect 184204 3606 184256 3612
rect 184860 3602 184888 57462
rect 185596 56710 185624 59758
rect 186424 57526 186452 59758
rect 187344 57798 187372 59758
rect 186964 57792 187016 57798
rect 186964 57734 187016 57740
rect 187332 57792 187384 57798
rect 187332 57734 187384 57740
rect 186412 57520 186464 57526
rect 186412 57462 186464 57468
rect 185584 56704 185636 56710
rect 185584 56646 185636 56652
rect 186228 10872 186280 10878
rect 186228 10814 186280 10820
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 186136 3596 186188 3602
rect 186136 3538 186188 3544
rect 182376 598 182588 626
rect 182376 490 182404 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 462 182404 490
rect 182560 480 182588 598
rect 183756 480 183784 3538
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 184952 480 184980 3334
rect 186148 480 186176 3538
rect 186240 3398 186268 10814
rect 186228 3392 186280 3398
rect 186228 3334 186280 3340
rect 186976 3126 187004 57734
rect 187608 57520 187660 57526
rect 187608 57462 187660 57468
rect 187620 3942 187648 57462
rect 188264 57458 188292 59758
rect 188252 57452 188304 57458
rect 188252 57394 188304 57400
rect 188344 57384 188396 57390
rect 188344 57326 188396 57332
rect 187608 3936 187660 3942
rect 187608 3878 187660 3884
rect 188356 3738 188384 57326
rect 189184 57118 189212 59758
rect 189172 57112 189224 57118
rect 189172 57054 189224 57060
rect 190276 57112 190328 57118
rect 190276 57054 190328 57060
rect 188988 10940 189040 10946
rect 188988 10882 189040 10888
rect 188344 3732 188396 3738
rect 188344 3674 188396 3680
rect 187332 3664 187384 3670
rect 187332 3606 187384 3612
rect 186964 3120 187016 3126
rect 186964 3062 187016 3068
rect 187344 480 187372 3606
rect 189000 3398 189028 10882
rect 190288 3874 190316 57054
rect 190276 3868 190328 3874
rect 190276 3810 190328 3816
rect 190380 3806 190408 59758
rect 191024 57526 191052 59758
rect 191944 57526 191972 59758
rect 191012 57520 191064 57526
rect 191012 57462 191064 57468
rect 191748 57520 191800 57526
rect 191748 57462 191800 57468
rect 191932 57520 191984 57526
rect 191932 57462 191984 57468
rect 193036 57520 193088 57526
rect 193036 57462 193088 57468
rect 191104 56704 191156 56710
rect 191104 56646 191156 56652
rect 190828 6656 190880 6662
rect 190828 6598 190880 6604
rect 190368 3800 190420 3806
rect 190368 3742 190420 3748
rect 188528 3392 188580 3398
rect 188528 3334 188580 3340
rect 188988 3392 189040 3398
rect 188988 3334 189040 3340
rect 188540 480 188568 3334
rect 189724 3120 189776 3126
rect 189724 3062 189776 3068
rect 189736 480 189764 3062
rect 190840 480 190868 6598
rect 191116 3398 191144 56646
rect 191760 3738 191788 57462
rect 192944 11008 192996 11014
rect 192944 10950 192996 10956
rect 191748 3732 191800 3738
rect 191748 3674 191800 3680
rect 191104 3392 191156 3398
rect 191104 3334 191156 3340
rect 192956 3330 192984 10950
rect 193048 4282 193076 57462
rect 193140 4350 193168 59758
rect 193692 57526 193720 59758
rect 194612 57526 194640 59758
rect 193680 57520 193732 57526
rect 193680 57462 193732 57468
rect 194508 57520 194560 57526
rect 194508 57462 194560 57468
rect 194600 57520 194652 57526
rect 194600 57462 194652 57468
rect 194416 9104 194468 9110
rect 194416 9046 194468 9052
rect 193128 4344 193180 4350
rect 193128 4286 193180 4292
rect 193036 4276 193088 4282
rect 193036 4218 193088 4224
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 192024 3324 192076 3330
rect 192024 3266 192076 3272
rect 192944 3324 192996 3330
rect 192944 3266 192996 3272
rect 192036 480 192064 3266
rect 193232 480 193260 3334
rect 194428 480 194456 9046
rect 194520 4418 194548 57462
rect 195612 10260 195664 10266
rect 195612 10202 195664 10208
rect 194508 4412 194560 4418
rect 194508 4354 194560 4360
rect 195624 480 195652 10202
rect 195808 4554 195836 59758
rect 196452 57526 196480 59758
rect 197372 57526 197400 59758
rect 195888 57520 195940 57526
rect 195888 57462 195940 57468
rect 196440 57520 196492 57526
rect 196440 57462 196492 57468
rect 197268 57520 197320 57526
rect 197268 57462 197320 57468
rect 197360 57520 197412 57526
rect 197360 57462 197412 57468
rect 195796 4548 195848 4554
rect 195796 4490 195848 4496
rect 195900 4486 195928 57462
rect 196624 57112 196676 57118
rect 196624 57054 196676 57060
rect 195888 4480 195940 4486
rect 195888 4422 195940 4428
rect 196636 4010 196664 57054
rect 197280 4622 197308 57462
rect 197912 9172 197964 9178
rect 197912 9114 197964 9120
rect 197268 4616 197320 4622
rect 197268 4558 197320 4564
rect 196624 4004 196676 4010
rect 196624 3946 196676 3952
rect 196808 3936 196860 3942
rect 196808 3878 196860 3884
rect 196820 480 196848 3878
rect 197924 480 197952 9114
rect 198568 4758 198596 59758
rect 199212 57526 199240 59758
rect 200132 57798 200160 59758
rect 200120 57792 200172 57798
rect 200120 57734 200172 57740
rect 200960 57526 200988 59758
rect 201316 57792 201368 57798
rect 201316 57734 201368 57740
rect 198648 57520 198700 57526
rect 198648 57462 198700 57468
rect 199200 57520 199252 57526
rect 199200 57462 199252 57468
rect 200028 57520 200080 57526
rect 200028 57462 200080 57468
rect 200948 57520 201000 57526
rect 200948 57462 201000 57468
rect 198556 4752 198608 4758
rect 198556 4694 198608 4700
rect 198660 4690 198688 57462
rect 199936 10192 199988 10198
rect 199936 10134 199988 10140
rect 198648 4684 198700 4690
rect 198648 4626 198700 4632
rect 199948 3398 199976 10134
rect 200040 5506 200068 57462
rect 200120 57452 200172 57458
rect 200120 57394 200172 57400
rect 200132 16574 200160 57394
rect 200132 16546 200344 16574
rect 200028 5500 200080 5506
rect 200028 5442 200080 5448
rect 199108 3392 199160 3398
rect 199108 3334 199160 3340
rect 199936 3392 199988 3398
rect 199936 3334 199988 3340
rect 199120 480 199148 3334
rect 200316 480 200344 16546
rect 201328 5438 201356 57734
rect 201880 57526 201908 59758
rect 202708 59758 202792 59786
rect 203684 59786 203712 60044
rect 204604 59786 204632 60044
rect 205524 59786 205552 60044
rect 203684 59758 203748 59786
rect 204604 59758 204668 59786
rect 201408 57520 201460 57526
rect 201408 57462 201460 57468
rect 201868 57520 201920 57526
rect 201868 57462 201920 57468
rect 201316 5432 201368 5438
rect 201316 5374 201368 5380
rect 201420 5370 201448 57462
rect 202604 10124 202656 10130
rect 202604 10066 202656 10072
rect 201500 9240 201552 9246
rect 201500 9182 201552 9188
rect 201408 5364 201460 5370
rect 201408 5306 201460 5312
rect 201512 480 201540 9182
rect 202616 3482 202644 10066
rect 202708 5234 202736 59758
rect 203720 57526 203748 59758
rect 204640 57526 204668 59758
rect 205468 59758 205552 59786
rect 206444 59786 206472 60044
rect 207364 59786 207392 60044
rect 208192 59786 208220 60044
rect 209112 59786 209140 60044
rect 210032 59786 210060 60044
rect 210952 59786 210980 60044
rect 211872 59786 211900 60044
rect 212792 59786 212820 60044
rect 213712 59786 213740 60044
rect 214632 59786 214660 60044
rect 215460 59786 215488 60044
rect 216380 59786 216408 60044
rect 217300 59786 217328 60044
rect 218220 59786 218248 60044
rect 219140 59786 219168 60044
rect 220060 59786 220088 60044
rect 220980 59786 221008 60044
rect 221900 59786 221928 60044
rect 222728 59786 222756 60044
rect 223648 59786 223676 60044
rect 224568 59786 224596 60044
rect 225488 59786 225516 60044
rect 226408 59786 226436 60044
rect 227328 59786 227356 60044
rect 228248 59786 228276 60044
rect 229168 59786 229196 60044
rect 229996 59786 230024 60044
rect 230916 59786 230944 60044
rect 231836 59786 231864 60044
rect 232756 59786 232784 60044
rect 233676 59786 233704 60044
rect 234596 59786 234624 60044
rect 235516 59786 235544 60044
rect 236436 59786 236464 60044
rect 237264 59786 237292 60044
rect 238184 59786 238212 60044
rect 239104 59786 239132 60044
rect 240024 59786 240052 60044
rect 240944 59786 240972 60044
rect 241864 59786 241892 60044
rect 242784 59786 242812 60044
rect 243704 59786 243732 60044
rect 244532 59786 244560 60044
rect 245452 59786 245480 60044
rect 246372 59786 246400 60044
rect 247292 59786 247320 60044
rect 248212 59786 248240 60044
rect 249132 59786 249160 60044
rect 250052 59786 250080 60044
rect 250972 59786 251000 60044
rect 251800 59786 251828 60044
rect 252720 59786 252748 60044
rect 253640 59786 253668 60044
rect 254560 59786 254588 60044
rect 255480 59786 255508 60044
rect 256400 59786 256428 60044
rect 257320 59786 257348 60044
rect 258240 59786 258268 60044
rect 259068 59786 259096 60044
rect 259988 59786 260016 60044
rect 260908 59786 260936 60044
rect 261828 59786 261856 60044
rect 262748 59786 262776 60044
rect 263668 59786 263696 60044
rect 264588 59786 264616 60044
rect 265508 59786 265536 60044
rect 266336 59786 266364 60044
rect 267256 59786 267284 60044
rect 268176 59786 268204 60044
rect 269096 59786 269124 60044
rect 270016 59786 270044 60044
rect 270936 59786 270964 60044
rect 271856 59786 271884 60044
rect 272776 59786 272804 60044
rect 273604 59786 273632 60044
rect 274524 59786 274552 60044
rect 206444 59758 206508 59786
rect 207364 59758 207428 59786
rect 208192 59758 208348 59786
rect 209112 59758 209176 59786
rect 210032 59758 210096 59786
rect 210952 59758 211016 59786
rect 211872 59758 211936 59786
rect 212792 59758 212856 59786
rect 213712 59758 213868 59786
rect 214632 59758 214696 59786
rect 215460 59758 215524 59786
rect 216380 59758 216628 59786
rect 217300 59758 217364 59786
rect 218220 59758 218284 59786
rect 219140 59758 219204 59786
rect 220060 59758 220124 59786
rect 220980 59758 221044 59786
rect 221900 59758 221964 59786
rect 222728 59758 222792 59786
rect 223648 59758 223712 59786
rect 224568 59758 224816 59786
rect 225488 59758 225552 59786
rect 226408 59758 226472 59786
rect 227328 59758 227668 59786
rect 228248 59758 228312 59786
rect 229168 59758 229232 59786
rect 229996 59758 230428 59786
rect 230916 59758 230980 59786
rect 231836 59758 231900 59786
rect 232756 59758 233188 59786
rect 233676 59758 233740 59786
rect 234596 59758 234660 59786
rect 235516 59758 235948 59786
rect 236436 59758 236500 59786
rect 237264 59758 237328 59786
rect 238184 59758 238248 59786
rect 239104 59758 239168 59786
rect 240024 59758 240088 59786
rect 240944 59758 241008 59786
rect 241864 59758 241928 59786
rect 242784 59758 242848 59786
rect 243704 59758 243768 59786
rect 244532 59758 244596 59786
rect 245452 59758 245516 59786
rect 246372 59758 246436 59786
rect 247292 59758 247356 59786
rect 248212 59758 248368 59786
rect 249132 59758 249196 59786
rect 250052 59758 250116 59786
rect 250972 59758 251128 59786
rect 251800 59758 251864 59786
rect 252720 59758 252784 59786
rect 253640 59758 253796 59786
rect 254560 59758 254624 59786
rect 255480 59758 255544 59786
rect 256400 59758 256648 59786
rect 257320 59758 257384 59786
rect 258240 59758 258304 59786
rect 259068 59758 259132 59786
rect 259988 59758 260052 59786
rect 260908 59758 260972 59786
rect 261828 59758 261892 59786
rect 262748 59758 262812 59786
rect 263668 59758 263732 59786
rect 264588 59758 264652 59786
rect 265508 59758 265572 59786
rect 266336 59758 266400 59786
rect 267256 59758 267688 59786
rect 268176 59758 268240 59786
rect 269096 59758 269160 59786
rect 270016 59758 270448 59786
rect 270936 59758 271000 59786
rect 271856 59758 271920 59786
rect 272776 59758 273116 59786
rect 273604 59758 273668 59786
rect 202788 57520 202840 57526
rect 202788 57462 202840 57468
rect 203708 57520 203760 57526
rect 203708 57462 203760 57468
rect 204168 57520 204220 57526
rect 204168 57462 204220 57468
rect 204628 57520 204680 57526
rect 204628 57462 204680 57468
rect 202800 5302 202828 57462
rect 202788 5296 202840 5302
rect 202788 5238 202840 5244
rect 202696 5228 202748 5234
rect 202696 5170 202748 5176
rect 204180 5166 204208 57462
rect 205088 9308 205140 9314
rect 205088 9250 205140 9256
rect 204168 5160 204220 5166
rect 204168 5102 204220 5108
rect 203892 4004 203944 4010
rect 203892 3946 203944 3952
rect 202616 3454 202736 3482
rect 202708 480 202736 3454
rect 203904 480 203932 3946
rect 205100 480 205128 9250
rect 205468 5030 205496 59758
rect 206480 57526 206508 59758
rect 205548 57520 205600 57526
rect 205548 57462 205600 57468
rect 206468 57520 206520 57526
rect 206468 57462 206520 57468
rect 206928 57520 206980 57526
rect 206928 57462 206980 57468
rect 205560 5098 205588 57462
rect 206836 10056 206888 10062
rect 206836 9998 206888 10004
rect 205548 5092 205600 5098
rect 205548 5034 205600 5040
rect 205456 5024 205508 5030
rect 205456 4966 205508 4972
rect 206848 3398 206876 9998
rect 206940 4962 206968 57462
rect 207400 57050 207428 59758
rect 207388 57044 207440 57050
rect 207388 56986 207440 56992
rect 208216 57044 208268 57050
rect 208216 56986 208268 56992
rect 206928 4956 206980 4962
rect 206928 4898 206980 4904
rect 208228 4894 208256 56986
rect 208216 4888 208268 4894
rect 208216 4830 208268 4836
rect 208320 4826 208348 59758
rect 209148 57526 209176 59758
rect 209136 57520 209188 57526
rect 209136 57462 209188 57468
rect 209688 57520 209740 57526
rect 209688 57462 209740 57468
rect 208584 9376 208636 9382
rect 208584 9318 208636 9324
rect 208308 4820 208360 4826
rect 208308 4762 208360 4768
rect 207388 3868 207440 3874
rect 207388 3810 207440 3816
rect 206192 3392 206244 3398
rect 206192 3334 206244 3340
rect 206836 3392 206888 3398
rect 206836 3334 206888 3340
rect 206204 480 206232 3334
rect 207400 480 207428 3810
rect 208596 480 208624 9318
rect 209700 6798 209728 57462
rect 210068 57050 210096 59758
rect 210988 57118 211016 59758
rect 211908 57458 211936 59758
rect 212828 57526 212856 59758
rect 212816 57520 212868 57526
rect 212816 57462 212868 57468
rect 213736 57520 213788 57526
rect 213736 57462 213788 57468
rect 211896 57452 211948 57458
rect 211896 57394 211948 57400
rect 210976 57112 211028 57118
rect 210976 57054 211028 57060
rect 210056 57044 210108 57050
rect 210056 56986 210108 56992
rect 213748 17406 213776 57462
rect 213736 17400 213788 17406
rect 213736 17342 213788 17348
rect 213840 12034 213868 59758
rect 214668 57526 214696 59758
rect 215496 57526 215524 59758
rect 214656 57520 214708 57526
rect 214656 57462 214708 57468
rect 215208 57520 215260 57526
rect 215208 57462 215260 57468
rect 215484 57520 215536 57526
rect 215484 57462 215536 57468
rect 216496 57520 216548 57526
rect 216496 57462 216548 57468
rect 214564 57044 214616 57050
rect 214564 56986 214616 56992
rect 214576 19990 214604 56986
rect 214564 19984 214616 19990
rect 214564 19926 214616 19932
rect 214564 17536 214616 17542
rect 214564 17478 214616 17484
rect 213828 12028 213880 12034
rect 213828 11970 213880 11976
rect 211068 9988 211120 9994
rect 211068 9930 211120 9936
rect 209688 6792 209740 6798
rect 209688 6734 209740 6740
rect 210976 3800 211028 3806
rect 210976 3742 211028 3748
rect 209780 3392 209832 3398
rect 209780 3334 209832 3340
rect 209792 480 209820 3334
rect 210988 480 211016 3742
rect 211080 3398 211108 9930
rect 213828 9920 213880 9926
rect 213828 9862 213880 9868
rect 212172 9444 212224 9450
rect 212172 9386 212224 9392
rect 211068 3392 211120 3398
rect 211068 3334 211120 3340
rect 212184 480 212212 9386
rect 213840 3398 213868 9862
rect 214472 3732 214524 3738
rect 214472 3674 214524 3680
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 213380 480 213408 3334
rect 214484 480 214512 3674
rect 214576 3670 214604 17478
rect 215220 12374 215248 57462
rect 215208 12368 215260 12374
rect 215208 12310 215260 12316
rect 216508 12306 216536 57462
rect 216496 12300 216548 12306
rect 216496 12242 216548 12248
rect 216600 12238 216628 59758
rect 217336 57526 217364 59758
rect 218256 57798 218284 59758
rect 218244 57792 218296 57798
rect 218244 57734 218296 57740
rect 217324 57520 217376 57526
rect 217324 57462 217376 57468
rect 217968 57520 218020 57526
rect 217968 57462 218020 57468
rect 217980 13598 218008 57462
rect 219176 57458 219204 59758
rect 220096 57526 220124 59758
rect 219992 57520 220044 57526
rect 219992 57462 220044 57468
rect 220084 57520 220136 57526
rect 220084 57462 220136 57468
rect 220728 57520 220780 57526
rect 220728 57462 220780 57468
rect 219164 57452 219216 57458
rect 219164 57394 219216 57400
rect 220004 55214 220032 57462
rect 220004 55186 220124 55214
rect 217968 13592 218020 13598
rect 217968 13534 218020 13540
rect 216588 12232 216640 12238
rect 216588 12174 216640 12180
rect 217968 9852 218020 9858
rect 217968 9794 218020 9800
rect 215668 9512 215720 9518
rect 215668 9454 215720 9460
rect 214564 3664 214616 3670
rect 214564 3606 214616 3612
rect 215680 480 215708 9454
rect 217980 3398 218008 9794
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 218060 4276 218112 4282
rect 218060 4218 218112 4224
rect 216864 3392 216916 3398
rect 216864 3334 216916 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 216876 480 216904 3334
rect 218072 480 218100 4218
rect 219268 480 219296 9522
rect 220096 6730 220124 55186
rect 220740 13462 220768 57462
rect 221016 56642 221044 59758
rect 221936 57458 221964 59758
rect 222764 57526 222792 59758
rect 222844 57792 222896 57798
rect 222844 57734 222896 57740
rect 222752 57520 222804 57526
rect 222752 57462 222804 57468
rect 221924 57452 221976 57458
rect 221924 57394 221976 57400
rect 221004 56636 221056 56642
rect 221004 56578 221056 56584
rect 222856 21486 222884 57734
rect 223684 57526 223712 59758
rect 223396 57520 223448 57526
rect 223396 57462 223448 57468
rect 223672 57520 223724 57526
rect 223672 57462 223724 57468
rect 223408 55214 223436 57462
rect 223408 55186 223528 55214
rect 222844 21480 222896 21486
rect 222844 21422 222896 21428
rect 220728 13456 220780 13462
rect 220728 13398 220780 13404
rect 223500 12170 223528 55186
rect 224788 22778 224816 59758
rect 225524 57798 225552 59758
rect 225512 57792 225564 57798
rect 225512 57734 225564 57740
rect 224868 57520 224920 57526
rect 224868 57462 224920 57468
rect 224776 22772 224828 22778
rect 224776 22714 224828 22720
rect 224224 16176 224276 16182
rect 224224 16118 224276 16124
rect 223488 12164 223540 12170
rect 223488 12106 223540 12112
rect 222752 9648 222804 9654
rect 222752 9590 222804 9596
rect 220084 6724 220136 6730
rect 220084 6666 220136 6672
rect 221556 4344 221608 4350
rect 221556 4286 221608 4292
rect 220452 3664 220504 3670
rect 220452 3606 220504 3612
rect 220464 480 220492 3606
rect 221568 480 221596 4286
rect 222764 480 222792 9590
rect 224236 3602 224264 16118
rect 224880 13530 224908 57462
rect 226444 54670 226472 59758
rect 226432 54664 226484 54670
rect 226432 54606 226484 54612
rect 227536 32428 227588 32434
rect 227536 32370 227588 32376
rect 224868 13524 224920 13530
rect 224868 13466 224920 13472
rect 226340 8900 226392 8906
rect 226340 8842 226392 8848
rect 225144 4412 225196 4418
rect 225144 4354 225196 4360
rect 224224 3596 224276 3602
rect 224224 3538 224276 3544
rect 223948 3324 224000 3330
rect 223948 3266 224000 3272
rect 223960 480 223988 3266
rect 225156 480 225184 4354
rect 226352 480 226380 8842
rect 227548 480 227576 32370
rect 227640 12102 227668 59758
rect 228284 56914 228312 59758
rect 229204 57526 229232 59758
rect 229192 57520 229244 57526
rect 229192 57462 229244 57468
rect 230296 57520 230348 57526
rect 230296 57462 230348 57468
rect 228364 57044 228416 57050
rect 228364 56986 228416 56992
rect 228272 56908 228324 56914
rect 228272 56850 228324 56856
rect 228376 13666 228404 56986
rect 229008 56908 229060 56914
rect 229008 56850 229060 56856
rect 228456 15972 228508 15978
rect 228456 15914 228508 15920
rect 228364 13660 228416 13666
rect 228364 13602 228416 13608
rect 227628 12096 227680 12102
rect 227628 12038 227680 12044
rect 228468 3330 228496 15914
rect 229020 14754 229048 56850
rect 229008 14748 229060 14754
rect 229008 14690 229060 14696
rect 229836 8832 229888 8838
rect 229836 8774 229888 8780
rect 228732 4480 228784 4486
rect 228732 4422 228784 4428
rect 228456 3324 228508 3330
rect 228456 3266 228508 3272
rect 228744 480 228772 4422
rect 229848 480 229876 8774
rect 230308 6526 230336 57462
rect 230296 6520 230348 6526
rect 230296 6462 230348 6468
rect 230400 6458 230428 59758
rect 230952 57526 230980 59758
rect 231872 57526 231900 59758
rect 230940 57520 230992 57526
rect 230940 57462 230992 57468
rect 231768 57520 231820 57526
rect 231768 57462 231820 57468
rect 231860 57520 231912 57526
rect 231860 57462 231912 57468
rect 233056 57520 233108 57526
rect 233056 57462 233108 57468
rect 231124 57452 231176 57458
rect 231124 57394 231176 57400
rect 231136 18698 231164 57394
rect 231124 18692 231176 18698
rect 231124 18634 231176 18640
rect 231676 18624 231728 18630
rect 231676 18566 231728 18572
rect 230388 6452 230440 6458
rect 230388 6394 230440 6400
rect 231688 3602 231716 18566
rect 231780 6390 231808 57462
rect 231768 6384 231820 6390
rect 231768 6326 231820 6332
rect 233068 6322 233096 57462
rect 233056 6316 233108 6322
rect 233056 6258 233108 6264
rect 233160 6254 233188 59758
rect 233712 57526 233740 59758
rect 234632 57798 234660 59758
rect 233884 57792 233936 57798
rect 233884 57734 233936 57740
rect 234620 57792 234672 57798
rect 234620 57734 234672 57740
rect 233700 57520 233752 57526
rect 233700 57462 233752 57468
rect 233896 50386 233924 57734
rect 234528 57520 234580 57526
rect 234528 57462 234580 57468
rect 233884 50380 233936 50386
rect 233884 50322 233936 50328
rect 233424 8764 233476 8770
rect 233424 8706 233476 8712
rect 233148 6248 233200 6254
rect 233148 6190 233200 6196
rect 232228 4548 232280 4554
rect 232228 4490 232280 4496
rect 231032 3596 231084 3602
rect 231032 3538 231084 3544
rect 231676 3596 231728 3602
rect 231676 3538 231728 3544
rect 231044 480 231072 3538
rect 232240 480 232268 4490
rect 233436 480 233464 8706
rect 234540 6186 234568 57462
rect 235920 14618 235948 59758
rect 236472 57458 236500 59758
rect 237300 57526 237328 59758
rect 237288 57520 237340 57526
rect 237288 57462 237340 57468
rect 238024 57520 238076 57526
rect 238024 57462 238076 57468
rect 236460 57452 236512 57458
rect 236460 57394 236512 57400
rect 238036 24138 238064 57462
rect 238220 57458 238248 59758
rect 238208 57452 238260 57458
rect 238208 57394 238260 57400
rect 238668 57452 238720 57458
rect 238668 57394 238720 57400
rect 238024 24132 238076 24138
rect 238024 24074 238076 24080
rect 238024 21412 238076 21418
rect 238024 21354 238076 21360
rect 235908 14612 235960 14618
rect 235908 14554 235960 14560
rect 237012 8696 237064 8702
rect 237012 8638 237064 8644
rect 234528 6180 234580 6186
rect 234528 6122 234580 6128
rect 235816 4616 235868 4622
rect 235816 4558 235868 4564
rect 234620 3596 234672 3602
rect 234620 3538 234672 3544
rect 234632 480 234660 3538
rect 235828 480 235856 4558
rect 237024 480 237052 8638
rect 238036 3670 238064 21354
rect 238680 13326 238708 57394
rect 239140 57050 239168 59758
rect 240060 57458 240088 59758
rect 240980 57458 241008 59758
rect 241900 57458 241928 59758
rect 240048 57452 240100 57458
rect 240048 57394 240100 57400
rect 240784 57452 240836 57458
rect 240784 57394 240836 57400
rect 240968 57452 241020 57458
rect 240968 57394 241020 57400
rect 241428 57452 241480 57458
rect 241428 57394 241480 57400
rect 241888 57452 241940 57458
rect 241888 57394 241940 57400
rect 242716 57452 242768 57458
rect 242716 57394 242768 57400
rect 239128 57044 239180 57050
rect 239128 56986 239180 56992
rect 240796 31074 240824 57394
rect 240784 31068 240836 31074
rect 240784 31010 240836 31016
rect 238668 13320 238720 13326
rect 238668 13262 238720 13268
rect 241440 11966 241468 57394
rect 242728 14686 242756 57394
rect 242716 14680 242768 14686
rect 242716 14622 242768 14628
rect 242716 14544 242768 14550
rect 242716 14486 242768 14492
rect 241428 11960 241480 11966
rect 241428 11902 241480 11908
rect 240508 8628 240560 8634
rect 240508 8570 240560 8576
rect 239312 4684 239364 4690
rect 239312 4626 239364 4632
rect 238116 3732 238168 3738
rect 238116 3674 238168 3680
rect 238024 3664 238076 3670
rect 238024 3606 238076 3612
rect 238128 480 238156 3674
rect 239324 480 239352 4626
rect 240520 480 240548 8570
rect 242728 3398 242756 14486
rect 242820 7138 242848 59758
rect 243740 57458 243768 59758
rect 244568 57458 244596 59758
rect 243728 57452 243780 57458
rect 243728 57394 243780 57400
rect 244188 57452 244240 57458
rect 244188 57394 244240 57400
rect 244556 57452 244608 57458
rect 244556 57394 244608 57400
rect 244096 8560 244148 8566
rect 244096 8502 244148 8508
rect 242808 7132 242860 7138
rect 242808 7074 242860 7080
rect 242900 4752 242952 4758
rect 242900 4694 242952 4700
rect 241704 3392 241756 3398
rect 241704 3334 241756 3340
rect 242716 3392 242768 3398
rect 242716 3334 242768 3340
rect 241716 480 241744 3334
rect 242912 480 242940 4694
rect 244108 480 244136 8502
rect 244200 7206 244228 57394
rect 245488 7342 245516 59758
rect 246408 57458 246436 59758
rect 247328 57458 247356 59758
rect 245568 57452 245620 57458
rect 245568 57394 245620 57400
rect 246396 57452 246448 57458
rect 246396 57394 246448 57400
rect 246948 57452 247000 57458
rect 246948 57394 247000 57400
rect 247316 57452 247368 57458
rect 247316 57394 247368 57400
rect 248236 57452 248288 57458
rect 248236 57394 248288 57400
rect 245476 7336 245528 7342
rect 245476 7278 245528 7284
rect 245580 7274 245608 57394
rect 246304 33788 246356 33794
rect 246304 33730 246356 33736
rect 245568 7268 245620 7274
rect 245568 7210 245620 7216
rect 244188 7200 244240 7206
rect 244188 7142 244240 7148
rect 246316 3398 246344 33730
rect 246960 7410 246988 57394
rect 247592 8492 247644 8498
rect 247592 8434 247644 8440
rect 246948 7404 247000 7410
rect 246948 7346 247000 7352
rect 246396 5500 246448 5506
rect 246396 5442 246448 5448
rect 245200 3392 245252 3398
rect 245200 3334 245252 3340
rect 246304 3392 246356 3398
rect 246304 3334 246356 3340
rect 245212 480 245240 3334
rect 246408 480 246436 5442
rect 247604 480 247632 8434
rect 248248 7478 248276 57394
rect 248340 7546 248368 59758
rect 249168 57050 249196 59758
rect 250088 57050 250116 59758
rect 249156 57044 249208 57050
rect 249156 56986 249208 56992
rect 249708 57044 249760 57050
rect 249708 56986 249760 56992
rect 250076 57044 250128 57050
rect 250076 56986 250128 56992
rect 250996 57044 251048 57050
rect 250996 56986 251048 56992
rect 249064 16040 249116 16046
rect 249064 15982 249116 15988
rect 248328 7540 248380 7546
rect 248328 7482 248380 7488
rect 248236 7472 248288 7478
rect 248236 7414 248288 7420
rect 248788 3936 248840 3942
rect 248788 3878 248840 3884
rect 248800 480 248828 3878
rect 249076 3738 249104 15982
rect 249720 8294 249748 56986
rect 249708 8288 249760 8294
rect 249708 8230 249760 8236
rect 251008 8226 251036 56986
rect 250996 8220 251048 8226
rect 250996 8162 251048 8168
rect 251100 8158 251128 59758
rect 251836 57050 251864 59758
rect 252756 57050 252784 59758
rect 251824 57044 251876 57050
rect 251824 56986 251876 56992
rect 252468 57044 252520 57050
rect 252468 56986 252520 56992
rect 252744 57044 252796 57050
rect 252744 56986 252796 56992
rect 251180 8424 251232 8430
rect 251180 8366 251232 8372
rect 251088 8152 251140 8158
rect 251088 8094 251140 8100
rect 249984 5432 250036 5438
rect 249984 5374 250036 5380
rect 249064 3732 249116 3738
rect 249064 3674 249116 3680
rect 249996 480 250024 5374
rect 251192 480 251220 8366
rect 252480 8090 252508 56986
rect 252468 8084 252520 8090
rect 252468 8026 252520 8032
rect 253768 7954 253796 59758
rect 254596 57050 254624 59758
rect 255516 57050 255544 59758
rect 253848 57044 253900 57050
rect 253848 56986 253900 56992
rect 254584 57044 254636 57050
rect 254584 56986 254636 56992
rect 255228 57044 255280 57050
rect 255228 56986 255280 56992
rect 255504 57044 255556 57050
rect 255504 56986 255556 56992
rect 256516 57044 256568 57050
rect 256516 56986 256568 56992
rect 253860 8022 253888 56986
rect 253848 8016 253900 8022
rect 253848 7958 253900 7964
rect 253756 7948 253808 7954
rect 253756 7890 253808 7896
rect 255240 7886 255268 56986
rect 255964 13728 256016 13734
rect 255964 13670 256016 13676
rect 255228 7880 255280 7886
rect 255228 7822 255280 7828
rect 253480 5364 253532 5370
rect 253480 5306 253532 5312
rect 252376 3800 252428 3806
rect 252376 3742 252428 3748
rect 252388 480 252416 3742
rect 253492 480 253520 5306
rect 255872 3732 255924 3738
rect 255872 3674 255924 3680
rect 254676 3392 254728 3398
rect 254676 3334 254728 3340
rect 254688 480 254716 3334
rect 255884 480 255912 3674
rect 255976 3398 256004 13670
rect 256528 7818 256556 56986
rect 256516 7812 256568 7818
rect 256516 7754 256568 7760
rect 256620 7750 256648 59758
rect 257356 57050 257384 59758
rect 258276 57118 258304 59758
rect 258264 57112 258316 57118
rect 258264 57054 258316 57060
rect 257344 57044 257396 57050
rect 257344 56986 257396 56992
rect 257988 57044 258040 57050
rect 257988 56986 258040 56992
rect 256608 7744 256660 7750
rect 256608 7686 256660 7692
rect 258000 7682 258028 56986
rect 259104 56982 259132 59758
rect 260024 57118 260052 59758
rect 259368 57112 259420 57118
rect 259368 57054 259420 57060
rect 260012 57112 260064 57118
rect 260012 57054 260064 57060
rect 260748 57112 260800 57118
rect 260748 57054 260800 57060
rect 259092 56976 259144 56982
rect 259092 56918 259144 56924
rect 259276 14952 259328 14958
rect 259276 14894 259328 14900
rect 257988 7676 258040 7682
rect 257988 7618 258040 7624
rect 257068 5296 257120 5302
rect 257068 5238 257120 5244
rect 255964 3392 256016 3398
rect 255964 3334 256016 3340
rect 257080 480 257108 5238
rect 259288 3602 259316 14894
rect 259380 7614 259408 57054
rect 260104 37936 260156 37942
rect 260104 37878 260156 37884
rect 259368 7608 259420 7614
rect 259368 7550 259420 7556
rect 260116 3670 260144 37878
rect 260656 13252 260708 13258
rect 260656 13194 260708 13200
rect 260564 5228 260616 5234
rect 260564 5170 260616 5176
rect 260104 3664 260156 3670
rect 260104 3606 260156 3612
rect 258264 3596 258316 3602
rect 258264 3538 258316 3544
rect 259276 3596 259328 3602
rect 259276 3538 259328 3544
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 258276 480 258304 3538
rect 259472 480 259500 3538
rect 260576 2666 260604 5170
rect 260668 3602 260696 13194
rect 260760 11762 260788 57054
rect 260944 56778 260972 59758
rect 260932 56772 260984 56778
rect 260932 56714 260984 56720
rect 261864 56030 261892 59758
rect 262784 57118 262812 59758
rect 263704 57118 263732 59758
rect 262772 57112 262824 57118
rect 262772 57054 262824 57060
rect 263508 57112 263560 57118
rect 263508 57054 263560 57060
rect 263692 57112 263744 57118
rect 263692 57054 263744 57060
rect 262864 56364 262916 56370
rect 262864 56306 262916 56312
rect 261852 56024 261904 56030
rect 261852 55966 261904 55972
rect 260748 11756 260800 11762
rect 260748 11698 260800 11704
rect 262876 3602 262904 56306
rect 263520 13122 263548 57054
rect 264244 57044 264296 57050
rect 264244 56986 264296 56992
rect 263508 13116 263560 13122
rect 263508 13058 263560 13064
rect 264256 6050 264284 56986
rect 264624 56982 264652 59758
rect 264888 57112 264940 57118
rect 264888 57054 264940 57060
rect 264612 56976 264664 56982
rect 264612 56918 264664 56924
rect 264900 14482 264928 57054
rect 265544 55962 265572 59758
rect 266372 57118 266400 59758
rect 266360 57112 266412 57118
rect 266360 57054 266412 57060
rect 267556 57112 267608 57118
rect 267556 57054 267608 57060
rect 265532 55956 265584 55962
rect 265532 55898 265584 55904
rect 267004 16108 267056 16114
rect 267004 16050 267056 16056
rect 264888 14476 264940 14482
rect 264888 14418 264940 14424
rect 264244 6044 264296 6050
rect 264244 5986 264296 5992
rect 265348 5976 265400 5982
rect 265348 5918 265400 5924
rect 264152 5160 264204 5166
rect 264152 5102 264204 5108
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 261760 3596 261812 3602
rect 261760 3538 261812 3544
rect 262864 3596 262916 3602
rect 262864 3538 262916 3544
rect 260576 2638 260696 2666
rect 260668 480 260696 2638
rect 261772 480 261800 3538
rect 262968 480 262996 3606
rect 264164 480 264192 5102
rect 265360 480 265388 5918
rect 267016 3942 267044 16050
rect 267568 15910 267596 57054
rect 267556 15904 267608 15910
rect 267556 15846 267608 15852
rect 267660 4282 267688 59758
rect 268212 57118 268240 59758
rect 269132 57118 269160 59758
rect 268200 57112 268252 57118
rect 268200 57054 268252 57060
rect 269028 57112 269080 57118
rect 269028 57054 269080 57060
rect 269120 57112 269172 57118
rect 269120 57054 269172 57060
rect 270316 57112 270368 57118
rect 270316 57054 270368 57060
rect 268936 20052 268988 20058
rect 268936 19994 268988 20000
rect 268948 6914 268976 19994
rect 268856 6886 268976 6914
rect 267740 5092 267792 5098
rect 267740 5034 267792 5040
rect 267648 4276 267700 4282
rect 267648 4218 267700 4224
rect 267004 3936 267056 3942
rect 267004 3878 267056 3884
rect 266544 3800 266596 3806
rect 266544 3742 266596 3748
rect 266556 480 266584 3742
rect 267752 480 267780 5034
rect 268856 480 268884 6886
rect 269040 4350 269068 57054
rect 270328 4418 270356 57054
rect 270420 4486 270448 59758
rect 270972 57118 271000 59758
rect 271892 57118 271920 59758
rect 270960 57112 271012 57118
rect 270960 57054 271012 57060
rect 271788 57112 271840 57118
rect 271788 57054 271840 57060
rect 271880 57112 271932 57118
rect 271880 57054 271932 57060
rect 271144 26920 271196 26926
rect 271144 26862 271196 26868
rect 270408 4480 270460 4486
rect 270408 4422 270460 4428
rect 270316 4412 270368 4418
rect 270316 4354 270368 4360
rect 269028 4344 269080 4350
rect 269028 4286 269080 4292
rect 271156 3874 271184 26862
rect 271236 5024 271288 5030
rect 271236 4966 271288 4972
rect 271144 3868 271196 3874
rect 271144 3810 271196 3816
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 270052 480 270080 3334
rect 271248 480 271276 4966
rect 271800 4554 271828 57054
rect 272432 6112 272484 6118
rect 272432 6054 272484 6060
rect 271788 4548 271840 4554
rect 271788 4490 271840 4496
rect 272444 480 272472 6054
rect 273088 4690 273116 59758
rect 273640 57118 273668 59758
rect 274468 59758 274552 59786
rect 275444 59786 275472 60044
rect 276364 59786 276392 60044
rect 277284 59786 277312 60044
rect 275444 59758 275508 59786
rect 276364 59758 276428 59786
rect 273168 57112 273220 57118
rect 273168 57054 273220 57060
rect 273628 57112 273680 57118
rect 273628 57054 273680 57060
rect 273076 4684 273128 4690
rect 273076 4626 273128 4632
rect 273180 4622 273208 57054
rect 274364 14816 274416 14822
rect 274364 14758 274416 14764
rect 273168 4616 273220 4622
rect 273168 4558 273220 4564
rect 274376 3602 274404 14758
rect 274468 5506 274496 59758
rect 275480 57118 275508 59758
rect 276400 57118 276428 59758
rect 277228 59758 277312 59786
rect 278204 59786 278232 60044
rect 279124 59786 279152 60044
rect 280044 59786 280072 60044
rect 280964 59786 280992 60044
rect 281792 59786 281820 60044
rect 282712 59786 282740 60044
rect 283632 59786 283660 60044
rect 284552 59786 284580 60044
rect 285472 59786 285500 60044
rect 286392 59786 286420 60044
rect 287312 59786 287340 60044
rect 288232 59786 288260 60044
rect 289060 59786 289088 60044
rect 289980 59786 290008 60044
rect 290900 59786 290928 60044
rect 291820 59786 291848 60044
rect 292740 59786 292768 60044
rect 293660 59786 293688 60044
rect 294580 59786 294608 60044
rect 278204 59758 278268 59786
rect 279124 59758 279188 59786
rect 280044 59758 280108 59786
rect 280964 59758 281028 59786
rect 281792 59758 281856 59786
rect 282712 59758 282776 59786
rect 283632 59758 283696 59786
rect 274548 57112 274600 57118
rect 274548 57054 274600 57060
rect 275468 57112 275520 57118
rect 275468 57054 275520 57060
rect 275928 57112 275980 57118
rect 275928 57054 275980 57060
rect 276388 57112 276440 57118
rect 276388 57054 276440 57060
rect 274456 5500 274508 5506
rect 274456 5442 274508 5448
rect 274560 4758 274588 57054
rect 275940 5438 275968 57054
rect 277124 12436 277176 12442
rect 277124 12378 277176 12384
rect 275928 5432 275980 5438
rect 275928 5374 275980 5380
rect 274824 4956 274876 4962
rect 274824 4898 274876 4904
rect 274548 4752 274600 4758
rect 274548 4694 274600 4700
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 274364 3596 274416 3602
rect 274364 3538 274416 3544
rect 273640 480 273668 3538
rect 274836 480 274864 4898
rect 277136 3602 277164 12378
rect 277228 5302 277256 59758
rect 278240 57118 278268 59758
rect 279160 57118 279188 59758
rect 277308 57112 277360 57118
rect 277308 57054 277360 57060
rect 278228 57112 278280 57118
rect 278228 57054 278280 57060
rect 278688 57112 278740 57118
rect 278688 57054 278740 57060
rect 279148 57112 279200 57118
rect 279148 57054 279200 57060
rect 279976 57112 280028 57118
rect 279976 57054 280028 57060
rect 277320 5370 277348 57054
rect 278044 17264 278096 17270
rect 278044 17206 278096 17212
rect 277308 5364 277360 5370
rect 277308 5306 277360 5312
rect 277216 5296 277268 5302
rect 277216 5238 277268 5244
rect 277216 3936 277268 3942
rect 277216 3878 277268 3884
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 276032 480 276060 3538
rect 277228 1986 277256 3878
rect 278056 3602 278084 17206
rect 278700 5234 278728 57054
rect 279516 6860 279568 6866
rect 279516 6802 279568 6808
rect 278688 5228 278740 5234
rect 278688 5170 278740 5176
rect 278320 4888 278372 4894
rect 278320 4830 278372 4836
rect 278044 3596 278096 3602
rect 278044 3538 278096 3544
rect 277136 1958 277256 1986
rect 277136 480 277164 1958
rect 278332 480 278360 4830
rect 279528 480 279556 6802
rect 279988 5166 280016 57054
rect 279976 5160 280028 5166
rect 279976 5102 280028 5108
rect 280080 5098 280108 59758
rect 281000 57118 281028 59758
rect 281828 57118 281856 59758
rect 280988 57112 281040 57118
rect 280988 57054 281040 57060
rect 281448 57112 281500 57118
rect 281448 57054 281500 57060
rect 281816 57112 281868 57118
rect 281816 57054 281868 57060
rect 280804 56092 280856 56098
rect 280804 56034 280856 56040
rect 280068 5092 280120 5098
rect 280068 5034 280120 5040
rect 280816 3738 280844 56034
rect 281460 5030 281488 57054
rect 281448 5024 281500 5030
rect 281448 4966 281500 4972
rect 282748 4894 282776 59758
rect 283668 57118 283696 59758
rect 284312 59758 284580 59786
rect 284680 59758 285500 59786
rect 285692 59758 286420 59786
rect 287256 59758 287340 59786
rect 288176 59758 288260 59786
rect 289004 59758 289088 59786
rect 289924 59758 290008 59786
rect 290844 59758 290928 59786
rect 291764 59758 291848 59786
rect 292684 59758 292768 59786
rect 293604 59758 293688 59786
rect 294524 59758 294608 59786
rect 295340 59832 295392 59838
rect 295500 59786 295528 60044
rect 296328 59838 296356 60044
rect 295340 59774 295392 59780
rect 282828 57112 282880 57118
rect 282828 57054 282880 57060
rect 283656 57112 283708 57118
rect 283656 57054 283708 57060
rect 284208 57112 284260 57118
rect 284208 57054 284260 57060
rect 282840 4962 282868 57054
rect 284116 9784 284168 9790
rect 284116 9726 284168 9732
rect 282828 4956 282880 4962
rect 282828 4898 282880 4904
rect 282736 4888 282788 4894
rect 282736 4830 282788 4836
rect 281908 4820 281960 4826
rect 281908 4762 281960 4768
rect 280804 3732 280856 3738
rect 280804 3674 280856 3680
rect 280712 3596 280764 3602
rect 280712 3538 280764 3544
rect 280724 480 280752 3538
rect 281920 480 281948 4762
rect 284128 3262 284156 9726
rect 284220 4826 284248 57054
rect 284312 7070 284340 59758
rect 284680 45554 284708 59758
rect 284404 45526 284708 45554
rect 284404 8974 284432 45526
rect 285588 13388 285640 13394
rect 285588 13330 285640 13336
rect 284392 8968 284444 8974
rect 284392 8910 284444 8916
rect 284300 7064 284352 7070
rect 284300 7006 284352 7012
rect 285404 6792 285456 6798
rect 285404 6734 285456 6740
rect 284208 4820 284260 4826
rect 284208 4762 284260 4768
rect 283104 3256 283156 3262
rect 283104 3198 283156 3204
rect 284116 3256 284168 3262
rect 284116 3198 284168 3204
rect 283116 480 283144 3198
rect 284300 3052 284352 3058
rect 284300 2994 284352 3000
rect 284312 480 284340 2994
rect 285416 480 285444 6734
rect 285600 3058 285628 13330
rect 285692 9042 285720 59758
rect 287256 57186 287284 59758
rect 288176 57594 288204 59758
rect 289004 57662 289032 59758
rect 289924 57730 289952 59758
rect 290844 57866 290872 59758
rect 291764 57934 291792 59758
rect 291752 57928 291804 57934
rect 291752 57870 291804 57876
rect 290832 57860 290884 57866
rect 290832 57802 290884 57808
rect 289912 57724 289964 57730
rect 289912 57666 289964 57672
rect 288992 57656 289044 57662
rect 288992 57598 289044 57604
rect 288164 57588 288216 57594
rect 288164 57530 288216 57536
rect 288256 57588 288308 57594
rect 288256 57530 288308 57536
rect 287244 57180 287296 57186
rect 287244 57122 287296 57128
rect 286324 57112 286376 57118
rect 286324 57054 286376 57060
rect 285680 9036 285732 9042
rect 285680 8978 285732 8984
rect 286336 5982 286364 57054
rect 287796 57044 287848 57050
rect 287796 56986 287848 56992
rect 287704 56636 287756 56642
rect 287704 56578 287756 56584
rect 286600 6792 286652 6798
rect 286600 6734 286652 6740
rect 286324 5976 286376 5982
rect 286324 5918 286376 5924
rect 285588 3052 285640 3058
rect 285588 2994 285640 3000
rect 286612 480 286640 6734
rect 287716 6662 287744 56578
rect 287808 11898 287836 56986
rect 288268 56642 288296 57530
rect 292684 57050 292712 59758
rect 288440 57044 288492 57050
rect 288440 56986 288492 56992
rect 292672 57044 292724 57050
rect 292672 56986 292724 56992
rect 288256 56636 288308 56642
rect 288256 56578 288308 56584
rect 288452 54602 288480 56986
rect 291936 56976 291988 56982
rect 291936 56918 291988 56924
rect 289084 56908 289136 56914
rect 289084 56850 289136 56856
rect 288440 54596 288492 54602
rect 288440 54538 288492 54544
rect 288440 19984 288492 19990
rect 288440 19926 288492 19932
rect 288452 16574 288480 19926
rect 288452 16546 289032 16574
rect 287796 11892 287848 11898
rect 287796 11834 287848 11840
rect 287704 6656 287756 6662
rect 287704 6598 287756 6604
rect 287796 3732 287848 3738
rect 287796 3674 287848 3680
rect 287808 480 287836 3674
rect 289004 480 289032 16546
rect 289096 11830 289124 56850
rect 291844 56636 291896 56642
rect 291844 56578 291896 56584
rect 289084 11824 289136 11830
rect 289084 11766 289136 11772
rect 290188 6656 290240 6662
rect 290188 6598 290240 6604
rect 290200 480 290228 6598
rect 291856 6594 291884 56578
rect 291948 13190 291976 56918
rect 293604 56166 293632 59758
rect 294524 56234 294552 59758
rect 294512 56228 294564 56234
rect 294512 56170 294564 56176
rect 293592 56160 293644 56166
rect 293592 56102 293644 56108
rect 294604 29640 294656 29646
rect 294604 29582 294656 29588
rect 291936 13184 291988 13190
rect 291936 13126 291988 13132
rect 291844 6588 291896 6594
rect 291844 6530 291896 6536
rect 293684 6588 293736 6594
rect 293684 6530 293736 6536
rect 292580 6044 292632 6050
rect 292580 5986 292632 5992
rect 291384 3188 291436 3194
rect 291384 3130 291436 3136
rect 291396 480 291424 3130
rect 292592 480 292620 5986
rect 293696 480 293724 6530
rect 294616 3942 294644 29582
rect 295352 14890 295380 59774
rect 295444 59758 295528 59786
rect 296316 59832 296368 59838
rect 297248 59786 297276 60044
rect 296316 59774 296368 59780
rect 297192 59758 297276 59786
rect 298168 59786 298196 60044
rect 299088 59786 299116 60044
rect 300008 59786 300036 60044
rect 300928 59922 300956 60044
rect 298168 59758 298232 59786
rect 295444 25566 295472 59758
rect 297192 56642 297220 59758
rect 297180 56636 297232 56642
rect 297180 56578 297232 56584
rect 298100 55752 298152 55758
rect 298100 55694 298152 55700
rect 295432 25560 295484 25566
rect 295432 25502 295484 25508
rect 295984 25560 296036 25566
rect 295984 25502 296036 25508
rect 295340 14884 295392 14890
rect 295340 14826 295392 14832
rect 294604 3936 294656 3942
rect 294604 3878 294656 3884
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 294892 480 294920 3810
rect 295996 3806 296024 25502
rect 298112 16182 298140 55694
rect 298204 35222 298232 59758
rect 299032 59758 299116 59786
rect 299492 59758 300036 59786
rect 300872 59894 300956 59922
rect 299032 55758 299060 59758
rect 299020 55752 299072 55758
rect 299020 55694 299072 55700
rect 298192 35216 298244 35222
rect 298192 35158 298244 35164
rect 298744 35216 298796 35222
rect 298744 35158 298796 35164
rect 298100 16176 298152 16182
rect 298100 16118 298152 16124
rect 296076 6724 296128 6730
rect 296076 6666 296128 6672
rect 297272 6724 297324 6730
rect 297272 6666 297324 6672
rect 295984 3800 296036 3806
rect 295984 3742 296036 3748
rect 296088 480 296116 6666
rect 297284 480 297312 6666
rect 298468 3800 298520 3806
rect 298468 3742 298520 3748
rect 298480 480 298508 3742
rect 298756 3194 298784 35158
rect 299492 17542 299520 59758
rect 300872 57594 300900 59894
rect 301848 59786 301876 60044
rect 302768 59786 302796 60044
rect 300964 59758 301876 59786
rect 302344 59758 302796 59786
rect 303596 59786 303624 60044
rect 304516 59786 304544 60044
rect 305436 59786 305464 60044
rect 303596 59758 303660 59786
rect 300860 57588 300912 57594
rect 300860 57530 300912 57536
rect 299480 17536 299532 17542
rect 299480 17478 299532 17484
rect 299480 17400 299532 17406
rect 299480 17342 299532 17348
rect 298836 17332 298888 17338
rect 298836 17274 298888 17280
rect 298848 3670 298876 17274
rect 299492 16574 299520 17342
rect 299492 16546 299704 16574
rect 298836 3664 298888 3670
rect 298836 3606 298888 3612
rect 298744 3188 298796 3194
rect 298744 3130 298796 3136
rect 299676 480 299704 16546
rect 300964 9110 300992 59758
rect 302344 9178 302372 59758
rect 303160 12028 303212 12034
rect 303160 11970 303212 11976
rect 302332 9172 302384 9178
rect 302332 9114 302384 9120
rect 300952 9104 301004 9110
rect 300952 9046 301004 9052
rect 300768 6044 300820 6050
rect 300768 5986 300820 5992
rect 300780 480 300808 5986
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 301976 480 302004 3878
rect 303172 480 303200 11970
rect 303632 9246 303660 59758
rect 303724 59758 304544 59786
rect 305012 59758 305464 59786
rect 306356 59786 306384 60044
rect 307276 59786 307304 60044
rect 308196 59786 308224 60044
rect 306356 59758 306512 59786
rect 303724 9314 303752 59758
rect 305012 9382 305040 59758
rect 305644 57656 305696 57662
rect 305644 57598 305696 57604
rect 305000 9376 305052 9382
rect 305000 9318 305052 9324
rect 303712 9308 303764 9314
rect 303712 9250 303764 9256
rect 303620 9240 303672 9246
rect 303620 9182 303672 9188
rect 305656 6118 305684 57598
rect 306380 12368 306432 12374
rect 306380 12310 306432 12316
rect 306288 12028 306340 12034
rect 306288 11970 306340 11976
rect 305644 6112 305696 6118
rect 305644 6054 305696 6060
rect 304356 5976 304408 5982
rect 304356 5918 304408 5924
rect 304368 480 304396 5918
rect 306300 3398 306328 11970
rect 305552 3392 305604 3398
rect 305552 3334 305604 3340
rect 306288 3392 306340 3398
rect 306288 3334 306340 3340
rect 305564 480 305592 3334
rect 306392 490 306420 12310
rect 306484 9450 306512 59758
rect 306576 59758 307304 59786
rect 307772 59758 308224 59786
rect 309116 59786 309144 60044
rect 310036 59786 310064 60044
rect 310864 59786 310892 60044
rect 311784 59786 311812 60044
rect 312704 59786 312732 60044
rect 309116 59758 309364 59786
rect 306576 9518 306604 59758
rect 307772 9586 307800 59758
rect 309232 56772 309284 56778
rect 309232 56714 309284 56720
rect 307760 9580 307812 9586
rect 307760 9522 307812 9528
rect 306564 9512 306616 9518
rect 306564 9454 306616 9460
rect 306472 9444 306524 9450
rect 306472 9386 306524 9392
rect 309244 8906 309272 56714
rect 309336 9654 309364 59758
rect 309980 59758 310064 59786
rect 310532 59758 310892 59786
rect 310992 59758 311812 59786
rect 311912 59758 312732 59786
rect 313372 59832 313424 59838
rect 313624 59786 313652 60044
rect 314544 59838 314572 60044
rect 313372 59774 313424 59780
rect 309980 56778 310008 59758
rect 309968 56772 310020 56778
rect 309968 56714 310020 56720
rect 309784 12300 309836 12306
rect 309784 12242 309836 12248
rect 309324 9648 309376 9654
rect 309324 9590 309376 9596
rect 309232 8900 309284 8906
rect 309232 8842 309284 8848
rect 307944 6112 307996 6118
rect 307944 6054 307996 6060
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 6054
rect 309048 4004 309100 4010
rect 309048 3946 309100 3952
rect 309060 480 309088 3946
rect 309796 490 309824 12242
rect 310532 8838 310560 59758
rect 310992 45554 311020 59758
rect 310624 45526 311020 45554
rect 310520 8832 310572 8838
rect 310520 8774 310572 8780
rect 310624 8770 310652 45526
rect 310612 8764 310664 8770
rect 310612 8706 310664 8712
rect 311912 8702 311940 59758
rect 311900 8696 311952 8702
rect 311900 8638 311952 8644
rect 313384 8566 313412 59774
rect 313476 59758 313652 59786
rect 314532 59832 314584 59838
rect 315464 59786 315492 60044
rect 316384 59786 316412 60044
rect 317304 59786 317332 60044
rect 318132 59786 318160 60044
rect 319052 59786 319080 60044
rect 319972 59786 320000 60044
rect 320892 59786 320920 60044
rect 321812 59922 321840 60044
rect 314532 59774 314584 59780
rect 314672 59758 315492 59786
rect 316052 59758 316412 59786
rect 316604 59758 317332 59786
rect 317432 59758 318160 59786
rect 318996 59758 319080 59786
rect 319916 59758 320000 59786
rect 320284 59758 320920 59786
rect 321572 59894 321840 59922
rect 313476 8634 313504 59758
rect 313832 12232 313884 12238
rect 313832 12174 313884 12180
rect 313464 8628 313516 8634
rect 313464 8570 313516 8576
rect 313372 8560 313424 8566
rect 313372 8502 313424 8508
rect 311440 5908 311492 5914
rect 311440 5850 311492 5856
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 5850
rect 312636 3392 312688 3398
rect 312636 3334 312688 3340
rect 312648 480 312676 3334
rect 313844 480 313872 12174
rect 314672 8498 314700 59758
rect 314660 8492 314712 8498
rect 314660 8434 314712 8440
rect 316052 8430 316080 59758
rect 316604 45554 316632 59758
rect 316144 45526 316632 45554
rect 316144 13734 316172 45526
rect 317432 14958 317460 59758
rect 318996 56370 319024 59758
rect 319916 57118 319944 59758
rect 319904 57112 319956 57118
rect 319904 57054 319956 57060
rect 318984 56364 319036 56370
rect 318984 56306 319036 56312
rect 318064 56160 318116 56166
rect 318064 56102 318116 56108
rect 317420 14952 317472 14958
rect 317420 14894 317472 14900
rect 316132 13728 316184 13734
rect 316132 13670 316184 13676
rect 317328 13592 317380 13598
rect 317328 13534 317380 13540
rect 316040 8424 316092 8430
rect 316040 8366 316092 8372
rect 315028 5840 315080 5846
rect 315028 5782 315080 5788
rect 315040 480 315068 5782
rect 316224 3664 316276 3670
rect 316224 3606 316276 3612
rect 316236 480 316264 3606
rect 317340 480 317368 13534
rect 318076 3942 318104 56102
rect 320180 21480 320232 21486
rect 320180 21422 320232 21428
rect 320192 16574 320220 21422
rect 320284 20058 320312 59758
rect 321572 57662 321600 59894
rect 322732 59786 322760 60044
rect 323652 59786 323680 60044
rect 321664 59758 322760 59786
rect 322952 59758 323680 59786
rect 324320 59832 324372 59838
rect 324572 59786 324600 60044
rect 325400 59838 325428 60044
rect 324320 59774 324372 59780
rect 321560 57656 321612 57662
rect 321560 57598 321612 57604
rect 320824 57588 320876 57594
rect 320824 57530 320876 57536
rect 320272 20052 320324 20058
rect 320272 19994 320324 20000
rect 320192 16546 320496 16574
rect 318156 14884 318208 14890
rect 318156 14826 318208 14832
rect 318064 3936 318116 3942
rect 318064 3878 318116 3884
rect 318168 3602 318196 14826
rect 318524 5772 318576 5778
rect 318524 5714 318576 5720
rect 318156 3596 318208 3602
rect 318156 3538 318208 3544
rect 318536 480 318564 5714
rect 319720 4072 319772 4078
rect 319720 4014 319772 4020
rect 319732 480 319760 4014
rect 320468 490 320496 16546
rect 320836 3806 320864 57530
rect 321664 12442 321692 59758
rect 322204 56228 322256 56234
rect 322204 56170 322256 56176
rect 321652 12436 321704 12442
rect 321652 12378 321704 12384
rect 322112 5704 322164 5710
rect 322112 5646 322164 5652
rect 320824 3800 320876 3806
rect 320824 3742 320876 3748
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 5646
rect 322216 3738 322244 56170
rect 322952 6866 322980 59758
rect 323584 19984 323636 19990
rect 323584 19926 323636 19932
rect 322940 6860 322992 6866
rect 322940 6802 322992 6808
rect 323596 3874 323624 19926
rect 324332 6798 324360 59774
rect 324516 59758 324600 59786
rect 325388 59832 325440 59838
rect 326320 59786 326348 60044
rect 327240 59786 327268 60044
rect 328160 59786 328188 60044
rect 329080 59786 329108 60044
rect 330000 59786 330028 60044
rect 330920 59786 330948 60044
rect 331840 59786 331868 60044
rect 325388 59774 325440 59780
rect 325712 59758 326348 59786
rect 327184 59758 327268 59786
rect 327460 59758 328188 59786
rect 328472 59758 329108 59786
rect 329852 59758 330028 59786
rect 330680 59758 330948 59786
rect 331324 59758 331868 59786
rect 332668 59786 332696 60044
rect 333588 59786 333616 60044
rect 334508 59786 334536 60044
rect 332668 59758 332732 59786
rect 324412 13660 324464 13666
rect 324412 13602 324464 13608
rect 324320 6792 324372 6798
rect 324320 6734 324372 6740
rect 323584 3868 323636 3874
rect 323584 3810 323636 3816
rect 323308 3800 323360 3806
rect 323308 3742 323360 3748
rect 322204 3732 322256 3738
rect 322204 3674 322256 3680
rect 323320 480 323348 3742
rect 324424 480 324452 13602
rect 324516 9790 324544 59758
rect 324504 9784 324556 9790
rect 324504 9726 324556 9732
rect 325608 6792 325660 6798
rect 325608 6734 325660 6740
rect 325620 480 325648 6734
rect 325712 6662 325740 59758
rect 327080 13456 327132 13462
rect 327080 13398 327132 13404
rect 325700 6656 325752 6662
rect 325700 6598 325752 6604
rect 326804 3936 326856 3942
rect 326804 3878 326856 3884
rect 326816 480 326844 3878
rect 327092 3482 327120 13398
rect 327184 6594 327212 59758
rect 327460 45554 327488 59758
rect 327276 45526 327488 45554
rect 327276 6730 327304 45526
rect 327264 6724 327316 6730
rect 327264 6666 327316 6672
rect 327172 6588 327224 6594
rect 327172 6530 327224 6536
rect 328472 6050 328500 59758
rect 328460 6044 328512 6050
rect 328460 5986 328512 5992
rect 329852 5982 329880 59758
rect 330680 45554 330708 59758
rect 331220 56296 331272 56302
rect 331220 56238 331272 56244
rect 329944 45526 330708 45554
rect 329944 6118 329972 45526
rect 329932 6112 329984 6118
rect 329932 6054 329984 6060
rect 329840 5976 329892 5982
rect 329840 5918 329892 5924
rect 329196 5636 329248 5642
rect 329196 5578 329248 5584
rect 327092 3454 328040 3482
rect 328012 480 328040 3454
rect 329208 480 329236 5578
rect 330392 3732 330444 3738
rect 330392 3674 330444 3680
rect 330404 480 330432 3674
rect 331232 490 331260 56238
rect 331324 5914 331352 59758
rect 332600 57656 332652 57662
rect 332600 57598 332652 57604
rect 331312 5908 331364 5914
rect 331312 5850 331364 5856
rect 332612 5778 332640 57598
rect 332704 5846 332732 59758
rect 333532 59758 333616 59786
rect 333992 59758 334536 59786
rect 335428 59786 335456 60044
rect 336348 59786 336376 60044
rect 337268 59786 337296 60044
rect 338188 59786 338216 60044
rect 335428 59758 335492 59786
rect 333532 57662 333560 59758
rect 333520 57656 333572 57662
rect 333520 57598 333572 57604
rect 332692 5840 332744 5846
rect 332692 5782 332744 5788
rect 332600 5772 332652 5778
rect 332600 5714 332652 5720
rect 333992 5710 334020 59758
rect 335360 57656 335412 57662
rect 335360 57598 335412 57604
rect 334072 18692 334124 18698
rect 334072 18634 334124 18640
rect 334084 16574 334112 18634
rect 334084 16546 334664 16574
rect 333980 5704 334032 5710
rect 333980 5646 334032 5652
rect 332692 5568 332744 5574
rect 332692 5510 332744 5516
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 5510
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 333900 480 333928 3538
rect 334636 490 334664 16546
rect 334716 13456 334768 13462
rect 334716 13398 334768 13404
rect 334728 3602 334756 13398
rect 335372 5642 335400 57598
rect 335464 6798 335492 59758
rect 336292 59758 336376 59786
rect 336752 59758 337296 59786
rect 338132 59758 338216 59786
rect 339108 59786 339136 60044
rect 339936 59786 339964 60044
rect 340856 59786 340884 60044
rect 341776 59786 341804 60044
rect 342696 59786 342724 60044
rect 343616 59786 343644 60044
rect 344536 59786 344564 60044
rect 345456 59786 345484 60044
rect 346376 59786 346404 60044
rect 347204 59786 347232 60044
rect 348124 59786 348152 60044
rect 349044 59786 349072 60044
rect 349964 59786 349992 60044
rect 350884 59786 350912 60044
rect 351804 59786 351832 60044
rect 352724 59786 352752 60044
rect 353644 59786 353672 60044
rect 354472 59786 354500 60044
rect 355392 59786 355420 60044
rect 356312 59786 356340 60044
rect 357232 59786 357260 60044
rect 358152 59786 358180 60044
rect 359072 59786 359100 60044
rect 359992 59786 360020 60044
rect 360912 59786 360940 60044
rect 361740 59786 361768 60044
rect 362660 59786 362688 60044
rect 363580 59786 363608 60044
rect 364500 59786 364528 60044
rect 365420 59786 365448 60044
rect 366340 59786 366368 60044
rect 367260 59786 367288 60044
rect 368180 59786 368208 60044
rect 369008 59786 369036 60044
rect 369928 59786 369956 60044
rect 370848 59786 370876 60044
rect 371768 59786 371796 60044
rect 372688 59786 372716 60044
rect 373608 59786 373636 60044
rect 374528 59786 374556 60044
rect 375448 59786 375476 60044
rect 376276 59786 376304 60044
rect 377196 59786 377224 60044
rect 378116 59786 378144 60044
rect 379036 59786 379064 60044
rect 379956 59786 379984 60044
rect 380876 59786 380904 60044
rect 381796 59786 381824 60044
rect 382716 59786 382744 60044
rect 383636 59786 383664 60044
rect 384464 59786 384492 60044
rect 385384 59786 385412 60044
rect 386304 59786 386332 60044
rect 339108 59758 339448 59786
rect 339936 59758 340000 59786
rect 340856 59758 340920 59786
rect 341776 59758 342208 59786
rect 342696 59758 342760 59786
rect 343616 59758 343680 59786
rect 344536 59758 344876 59786
rect 345456 59758 345520 59786
rect 346376 59758 346440 59786
rect 347204 59758 347268 59786
rect 348124 59758 348188 59786
rect 349044 59758 349108 59786
rect 349964 59758 350028 59786
rect 350884 59758 350948 59786
rect 351804 59758 351868 59786
rect 352724 59758 352788 59786
rect 353644 59758 353708 59786
rect 354472 59758 354536 59786
rect 355392 59758 355456 59786
rect 356312 59758 356376 59786
rect 357232 59758 357388 59786
rect 358152 59758 358216 59786
rect 359072 59758 359136 59786
rect 359992 59758 360148 59786
rect 360912 59758 360976 59786
rect 361740 59758 361804 59786
rect 362660 59758 362908 59786
rect 363580 59758 363644 59786
rect 364500 59758 364564 59786
rect 365420 59758 365668 59786
rect 366340 59758 366404 59786
rect 367260 59758 367324 59786
rect 368180 59758 368336 59786
rect 369008 59758 369072 59786
rect 369928 59758 369992 59786
rect 370848 59758 371188 59786
rect 371768 59758 371832 59786
rect 372688 59758 372752 59786
rect 373608 59758 373948 59786
rect 374528 59758 374592 59786
rect 375448 59758 375512 59786
rect 376276 59758 376708 59786
rect 377196 59758 377260 59786
rect 378116 59758 378180 59786
rect 379036 59758 379468 59786
rect 379956 59758 380020 59786
rect 380876 59758 380940 59786
rect 381796 59758 382228 59786
rect 382716 59758 382780 59786
rect 383636 59758 383700 59786
rect 384464 59758 384528 59786
rect 385384 59758 385448 59786
rect 336292 57662 336320 59758
rect 336280 57656 336332 57662
rect 336280 57598 336332 57604
rect 335452 6792 335504 6798
rect 335452 6734 335504 6740
rect 336752 5642 336780 59758
rect 335360 5636 335412 5642
rect 335360 5578 335412 5584
rect 336740 5636 336792 5642
rect 336740 5578 336792 5584
rect 338132 5574 338160 59758
rect 338672 12164 338724 12170
rect 338672 12106 338724 12112
rect 336280 5568 336332 5574
rect 336280 5510 336332 5516
rect 338120 5568 338172 5574
rect 338120 5510 338172 5516
rect 334716 3596 334768 3602
rect 334716 3538 334768 3544
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 5510
rect 337476 3868 337528 3874
rect 337476 3810 337528 3816
rect 337488 480 337516 3810
rect 338684 480 338712 12106
rect 339420 5574 339448 59758
rect 339972 57662 340000 59758
rect 340892 57662 340920 59758
rect 339960 57656 340012 57662
rect 339960 57598 340012 57604
rect 340788 57656 340840 57662
rect 340788 57598 340840 57604
rect 340880 57656 340932 57662
rect 340880 57598 340932 57604
rect 342076 57656 342128 57662
rect 342076 57598 342128 57604
rect 340144 54596 340196 54602
rect 340144 54538 340196 54544
rect 339408 5568 339460 5574
rect 339408 5510 339460 5516
rect 339868 5568 339920 5574
rect 339868 5510 339920 5516
rect 339880 480 339908 5510
rect 340156 4010 340184 54538
rect 340800 5574 340828 57598
rect 340880 13524 340932 13530
rect 340880 13466 340932 13472
rect 340788 5568 340840 5574
rect 340788 5510 340840 5516
rect 340144 4004 340196 4010
rect 340144 3946 340196 3952
rect 340892 3602 340920 13466
rect 342088 5710 342116 57598
rect 342180 6662 342208 59758
rect 342732 57662 342760 59758
rect 343652 57662 343680 59758
rect 342720 57656 342772 57662
rect 342720 57598 342772 57604
rect 343548 57656 343600 57662
rect 343548 57598 343600 57604
rect 343640 57656 343692 57662
rect 343640 57598 343692 57604
rect 342904 36576 342956 36582
rect 342904 36518 342956 36524
rect 342168 6656 342220 6662
rect 342168 6598 342220 6604
rect 342076 5704 342128 5710
rect 342076 5646 342128 5652
rect 340972 4140 341024 4146
rect 340972 4082 341024 4088
rect 340880 3596 340932 3602
rect 340880 3538 340932 3544
rect 340984 480 341012 4082
rect 342168 3596 342220 3602
rect 342168 3538 342220 3544
rect 342180 480 342208 3538
rect 342916 3398 342944 36518
rect 343560 6594 343588 57598
rect 343548 6588 343600 6594
rect 343548 6530 343600 6536
rect 344848 5914 344876 59758
rect 345492 57662 345520 59758
rect 346412 57662 346440 59758
rect 344928 57656 344980 57662
rect 344928 57598 344980 57604
rect 345480 57656 345532 57662
rect 345480 57598 345532 57604
rect 346308 57656 346360 57662
rect 346308 57598 346360 57604
rect 346400 57656 346452 57662
rect 346400 57598 346452 57604
rect 344836 5908 344888 5914
rect 344836 5850 344888 5856
rect 344940 5778 344968 57598
rect 345020 22772 345072 22778
rect 345020 22714 345072 22720
rect 345032 16574 345060 22714
rect 345032 16546 345336 16574
rect 344928 5772 344980 5778
rect 344928 5714 344980 5720
rect 343364 5568 343416 5574
rect 343364 5510 343416 5516
rect 342904 3392 342956 3398
rect 342904 3334 342956 3340
rect 343376 480 343404 5510
rect 344560 4004 344612 4010
rect 344560 3946 344612 3952
rect 344572 480 344600 3946
rect 345308 490 345336 16546
rect 346320 5642 346348 57598
rect 347240 56778 347268 59758
rect 348160 57662 348188 59758
rect 347596 57656 347648 57662
rect 347596 57598 347648 57604
rect 348148 57656 348200 57662
rect 348148 57598 348200 57604
rect 348976 57656 349028 57662
rect 348976 57598 349028 57604
rect 347228 56772 347280 56778
rect 347228 56714 347280 56720
rect 347608 5846 347636 57598
rect 347688 56772 347740 56778
rect 347688 56714 347740 56720
rect 347700 5982 347728 56714
rect 348988 6050 349016 57598
rect 349080 6118 349108 59758
rect 350000 56778 350028 59758
rect 350920 57662 350948 59758
rect 350908 57656 350960 57662
rect 350908 57598 350960 57604
rect 351736 57656 351788 57662
rect 351736 57598 351788 57604
rect 349988 56772 350040 56778
rect 349988 56714 350040 56720
rect 350448 56772 350500 56778
rect 350448 56714 350500 56720
rect 349160 50380 349212 50386
rect 349160 50322 349212 50328
rect 349172 16574 349200 50322
rect 349172 16546 349292 16574
rect 349068 6112 349120 6118
rect 349068 6054 349120 6060
rect 348976 6044 349028 6050
rect 348976 5986 349028 5992
rect 347688 5976 347740 5982
rect 347688 5918 347740 5924
rect 347596 5840 347648 5846
rect 347596 5782 347648 5788
rect 346952 5704 347004 5710
rect 346952 5646 347004 5652
rect 346308 5636 346360 5642
rect 346308 5578 346360 5584
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 5646
rect 348056 3392 348108 3398
rect 348056 3334 348108 3340
rect 348068 480 348096 3334
rect 349264 480 349292 16546
rect 350460 6866 350488 56714
rect 350448 6860 350500 6866
rect 350448 6802 350500 6808
rect 351748 6798 351776 57598
rect 351736 6792 351788 6798
rect 351736 6734 351788 6740
rect 351840 6730 351868 59758
rect 352760 56778 352788 59758
rect 353680 57662 353708 59758
rect 353668 57656 353720 57662
rect 353668 57598 353720 57604
rect 352748 56772 352800 56778
rect 352748 56714 352800 56720
rect 353208 56772 353260 56778
rect 353208 56714 353260 56720
rect 351920 54664 351972 54670
rect 351920 54606 351972 54612
rect 351932 16574 351960 54606
rect 351932 16546 352880 16574
rect 351828 6724 351880 6730
rect 351828 6666 351880 6672
rect 350448 6656 350500 6662
rect 350448 6598 350500 6604
rect 350460 480 350488 6598
rect 351644 3596 351696 3602
rect 351644 3538 351696 3544
rect 351656 480 351684 3538
rect 352852 480 352880 16546
rect 353220 6662 353248 56714
rect 353208 6656 353260 6662
rect 353208 6598 353260 6604
rect 354036 6588 354088 6594
rect 354036 6530 354088 6536
rect 354048 480 354076 6530
rect 354508 5574 354536 59758
rect 355428 57662 355456 59758
rect 356348 57662 356376 59758
rect 354588 57656 354640 57662
rect 354588 57598 354640 57604
rect 355416 57656 355468 57662
rect 355416 57598 355468 57604
rect 355968 57656 356020 57662
rect 355968 57598 356020 57604
rect 356336 57656 356388 57662
rect 356336 57598 356388 57604
rect 357256 57656 357308 57662
rect 357256 57598 357308 57604
rect 354600 6594 354628 57598
rect 355980 7070 356008 57598
rect 357268 18766 357296 57598
rect 357256 18760 357308 18766
rect 357256 18702 357308 18708
rect 356704 18692 356756 18698
rect 356704 18634 356756 18640
rect 356336 12096 356388 12102
rect 356336 12038 356388 12044
rect 355968 7064 356020 7070
rect 355968 7006 356020 7012
rect 354588 6588 354640 6594
rect 354588 6530 354640 6536
rect 354496 5568 354548 5574
rect 354496 5510 354548 5516
rect 355230 3360 355286 3369
rect 355230 3295 355286 3304
rect 355244 480 355272 3295
rect 356348 480 356376 12038
rect 356716 4078 356744 18634
rect 357360 12306 357388 59758
rect 358188 57662 358216 59758
rect 359108 57662 359136 59758
rect 358176 57656 358228 57662
rect 358176 57598 358228 57604
rect 358728 57656 358780 57662
rect 358728 57598 358780 57604
rect 359096 57656 359148 57662
rect 359096 57598 359148 57604
rect 360016 57656 360068 57662
rect 360016 57598 360068 57604
rect 358084 22772 358136 22778
rect 358084 22714 358136 22720
rect 357348 12300 357400 12306
rect 357348 12242 357400 12248
rect 357532 5704 357584 5710
rect 357532 5646 357584 5652
rect 356704 4072 356756 4078
rect 356704 4014 356756 4020
rect 357544 480 357572 5646
rect 358096 3670 358124 22714
rect 358740 8430 358768 57598
rect 359464 14748 359516 14754
rect 359464 14690 359516 14696
rect 358728 8424 358780 8430
rect 358728 8366 358780 8372
rect 358084 3664 358136 3670
rect 358084 3606 358136 3612
rect 358726 3496 358782 3505
rect 358726 3431 358782 3440
rect 358740 480 358768 3431
rect 359476 490 359504 14690
rect 360028 8498 360056 57598
rect 360120 8566 360148 59758
rect 360948 57662 360976 59758
rect 360936 57656 360988 57662
rect 360936 57598 360988 57604
rect 361488 57656 361540 57662
rect 361488 57598 361540 57604
rect 360844 14748 360896 14754
rect 360844 14690 360896 14696
rect 360108 8560 360160 8566
rect 360108 8502 360160 8508
rect 360016 8492 360068 8498
rect 360016 8434 360068 8440
rect 360856 3806 360884 14690
rect 361500 8634 361528 57598
rect 361776 56778 361804 59758
rect 361764 56772 361816 56778
rect 361764 56714 361816 56720
rect 362776 56772 362828 56778
rect 362776 56714 362828 56720
rect 362788 8702 362816 56714
rect 362880 8770 362908 59758
rect 363616 57662 363644 59758
rect 364536 57662 364564 59758
rect 363604 57656 363656 57662
rect 363604 57598 363656 57604
rect 364248 57656 364300 57662
rect 364248 57598 364300 57604
rect 364524 57656 364576 57662
rect 364524 57598 364576 57604
rect 365536 57656 365588 57662
rect 365536 57598 365588 57604
rect 363604 56296 363656 56302
rect 363604 56238 363656 56244
rect 362868 8764 362920 8770
rect 362868 8706 362920 8712
rect 362776 8696 362828 8702
rect 362776 8638 362828 8644
rect 361488 8628 361540 8634
rect 361488 8570 361540 8576
rect 363512 6520 363564 6526
rect 363512 6462 363564 6468
rect 361120 5772 361172 5778
rect 361120 5714 361172 5720
rect 360844 3800 360896 3806
rect 360844 3742 360896 3748
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 5714
rect 362314 3632 362370 3641
rect 362314 3567 362370 3576
rect 362328 480 362356 3567
rect 363524 480 363552 6462
rect 363616 3942 363644 56238
rect 364260 8838 364288 57598
rect 365548 8906 365576 57598
rect 365640 9654 365668 59758
rect 366376 57662 366404 59758
rect 367296 57662 367324 59758
rect 366364 57656 366416 57662
rect 366364 57598 366416 57604
rect 367008 57656 367060 57662
rect 367008 57598 367060 57604
rect 367284 57656 367336 57662
rect 367284 57598 367336 57604
rect 365628 9648 365680 9654
rect 365628 9590 365680 9596
rect 367020 9586 367048 57598
rect 367008 9580 367060 9586
rect 367008 9522 367060 9528
rect 368308 9450 368336 59758
rect 369044 57662 369072 59758
rect 369964 57662 369992 59758
rect 368388 57656 368440 57662
rect 368388 57598 368440 57604
rect 369032 57656 369084 57662
rect 369032 57598 369084 57604
rect 369768 57656 369820 57662
rect 369768 57598 369820 57604
rect 369952 57656 370004 57662
rect 369952 57598 370004 57604
rect 371056 57656 371108 57662
rect 371056 57598 371108 57604
rect 368400 9518 368428 57598
rect 368388 9512 368440 9518
rect 368388 9454 368440 9460
rect 368296 9444 368348 9450
rect 368296 9386 368348 9392
rect 369780 9382 369808 57598
rect 369768 9376 369820 9382
rect 369768 9318 369820 9324
rect 371068 9314 371096 57598
rect 371056 9308 371108 9314
rect 371056 9250 371108 9256
rect 371160 9246 371188 59758
rect 371804 57662 371832 59758
rect 372724 57662 372752 59758
rect 371792 57656 371844 57662
rect 371792 57598 371844 57604
rect 372528 57656 372580 57662
rect 372528 57598 372580 57604
rect 372712 57656 372764 57662
rect 372712 57598 372764 57604
rect 373816 57656 373868 57662
rect 373816 57598 373868 57604
rect 371884 39364 371936 39370
rect 371884 39306 371936 39312
rect 371148 9240 371200 9246
rect 371148 9182 371200 9188
rect 365536 8900 365588 8906
rect 365536 8842 365588 8848
rect 364248 8832 364300 8838
rect 364248 8774 364300 8780
rect 367008 6452 367060 6458
rect 367008 6394 367060 6400
rect 364616 5840 364668 5846
rect 364616 5782 364668 5788
rect 363604 3936 363656 3942
rect 363604 3878 363656 3884
rect 364628 480 364656 5782
rect 365810 3768 365866 3777
rect 365810 3703 365866 3712
rect 365824 480 365852 3703
rect 367020 480 367048 6394
rect 370596 6384 370648 6390
rect 370596 6326 370648 6332
rect 368204 5908 368256 5914
rect 368204 5850 368256 5856
rect 368216 480 368244 5850
rect 369400 3664 369452 3670
rect 369400 3606 369452 3612
rect 369412 480 369440 3606
rect 370608 480 370636 6326
rect 371700 5976 371752 5982
rect 371700 5918 371752 5924
rect 371712 480 371740 5918
rect 371896 3738 371924 39306
rect 372540 9178 372568 57598
rect 372528 9172 372580 9178
rect 372528 9114 372580 9120
rect 373828 9110 373856 57598
rect 373816 9104 373868 9110
rect 373816 9046 373868 9052
rect 373920 9042 373948 59758
rect 374564 57662 374592 59758
rect 375484 57866 375512 59758
rect 375472 57860 375524 57866
rect 375472 57802 375524 57808
rect 374644 57792 374696 57798
rect 374644 57734 374696 57740
rect 374552 57656 374604 57662
rect 374552 57598 374604 57604
rect 373908 9036 373960 9042
rect 373908 8978 373960 8984
rect 374656 6322 374684 57734
rect 375288 57656 375340 57662
rect 375288 57598 375340 57604
rect 375300 8974 375328 57598
rect 376024 40724 376076 40730
rect 376024 40666 376076 40672
rect 375288 8968 375340 8974
rect 375288 8910 375340 8916
rect 374092 6316 374144 6322
rect 374092 6258 374144 6264
rect 374644 6316 374696 6322
rect 374644 6258 374696 6264
rect 371884 3732 371936 3738
rect 371884 3674 371936 3680
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 374104 480 374132 6258
rect 375288 6044 375340 6050
rect 375288 5986 375340 5992
rect 375300 480 375328 5986
rect 376036 3874 376064 40666
rect 376680 12238 376708 59758
rect 377232 57662 377260 59758
rect 377404 57724 377456 57730
rect 377404 57666 377456 57672
rect 377220 57656 377272 57662
rect 377220 57598 377272 57604
rect 376668 12232 376720 12238
rect 376668 12174 376720 12180
rect 377416 4146 377444 57666
rect 378152 57662 378180 59758
rect 378048 57656 378100 57662
rect 378048 57598 378100 57604
rect 378140 57656 378192 57662
rect 378140 57598 378192 57604
rect 379336 57656 379388 57662
rect 379336 57598 379388 57604
rect 378060 13530 378088 57598
rect 378784 17468 378836 17474
rect 378784 17410 378836 17416
rect 378048 13524 378100 13530
rect 378048 13466 378100 13472
rect 377680 6248 377732 6254
rect 377680 6190 377732 6196
rect 377404 4140 377456 4146
rect 377404 4082 377456 4088
rect 376024 3868 376076 3874
rect 376024 3810 376076 3816
rect 376484 3800 376536 3806
rect 376484 3742 376536 3748
rect 376496 480 376524 3742
rect 377692 480 377720 6190
rect 378796 3398 378824 17410
rect 379348 17406 379376 57598
rect 379336 17400 379388 17406
rect 379336 17342 379388 17348
rect 379440 12170 379468 59758
rect 379992 57662 380020 59758
rect 380912 57798 380940 59758
rect 380900 57792 380952 57798
rect 380900 57734 380952 57740
rect 379980 57656 380032 57662
rect 379980 57598 380032 57604
rect 379428 12164 379480 12170
rect 379428 12106 379480 12112
rect 382200 12102 382228 59758
rect 382752 57186 382780 59758
rect 383672 57934 383700 59758
rect 383660 57928 383712 57934
rect 383660 57870 383712 57876
rect 384500 57526 384528 59758
rect 384856 57928 384908 57934
rect 384856 57870 384908 57876
rect 384488 57520 384540 57526
rect 384488 57462 384540 57468
rect 382740 57180 382792 57186
rect 382740 57122 382792 57128
rect 383568 57180 383620 57186
rect 383568 57122 383620 57128
rect 382924 56364 382976 56370
rect 382924 56306 382976 56312
rect 382188 12096 382240 12102
rect 382188 12038 382240 12044
rect 382372 6860 382424 6866
rect 382372 6802 382424 6808
rect 381176 6180 381228 6186
rect 381176 6122 381228 6128
rect 378876 6112 378928 6118
rect 378876 6054 378928 6060
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 378888 480 378916 6054
rect 379980 3868 380032 3874
rect 379980 3810 380032 3816
rect 379992 480 380020 3810
rect 381188 480 381216 6122
rect 382384 480 382412 6802
rect 382936 4010 382964 56306
rect 383580 13598 383608 57122
rect 383568 13592 383620 13598
rect 383568 13534 383620 13540
rect 384764 6316 384816 6322
rect 384764 6258 384816 6264
rect 382924 4004 382976 4010
rect 382924 3946 382976 3952
rect 383568 3936 383620 3942
rect 383568 3878 383620 3884
rect 383580 480 383608 3878
rect 384776 480 384804 6258
rect 384868 6186 384896 57870
rect 385420 57526 385448 59758
rect 386248 59758 386332 59786
rect 387224 59786 387252 60044
rect 388144 59786 388172 60044
rect 389064 59786 389092 60044
rect 389984 59786 390012 60044
rect 390904 59786 390932 60044
rect 391732 59786 391760 60044
rect 392652 59786 392680 60044
rect 393572 59786 393600 60044
rect 394492 59786 394520 60044
rect 395412 59786 395440 60044
rect 396332 59786 396360 60044
rect 397252 59786 397280 60044
rect 398172 59786 398200 60044
rect 399000 59786 399028 60044
rect 399920 59786 399948 60044
rect 400840 59786 400868 60044
rect 401760 59786 401788 60044
rect 402680 59786 402708 60044
rect 403600 59786 403628 60044
rect 404520 59786 404548 60044
rect 405440 59786 405468 60044
rect 406268 59786 406296 60044
rect 407188 59786 407216 60044
rect 408108 59786 408136 60044
rect 409028 59786 409056 60044
rect 387224 59758 387288 59786
rect 388144 59758 388208 59786
rect 389064 59758 389128 59786
rect 389984 59758 390048 59786
rect 390904 59758 390968 59786
rect 391732 59758 391888 59786
rect 392652 59758 392716 59786
rect 393572 59758 393636 59786
rect 394492 59758 394648 59786
rect 395412 59758 395476 59786
rect 396332 59758 396396 59786
rect 397252 59758 397316 59786
rect 398172 59758 398236 59786
rect 399000 59758 399064 59786
rect 399920 59758 400076 59786
rect 384948 57520 385000 57526
rect 384948 57462 385000 57468
rect 385408 57520 385460 57526
rect 385408 57462 385460 57468
rect 384856 6180 384908 6186
rect 384856 6122 384908 6128
rect 384960 5710 384988 57462
rect 385960 6792 386012 6798
rect 385960 6734 386012 6740
rect 384948 5704 385000 5710
rect 384948 5646 385000 5652
rect 385972 480 386000 6734
rect 386248 5846 386276 59758
rect 387260 57526 387288 59758
rect 388180 57526 388208 59758
rect 386328 57520 386380 57526
rect 386328 57462 386380 57468
rect 387248 57520 387300 57526
rect 387248 57462 387300 57468
rect 387708 57520 387760 57526
rect 387708 57462 387760 57468
rect 388168 57520 388220 57526
rect 388168 57462 388220 57468
rect 388996 57520 389048 57526
rect 388996 57462 389048 57468
rect 386236 5840 386288 5846
rect 386236 5782 386288 5788
rect 386340 5778 386368 57462
rect 387720 5914 387748 57462
rect 387800 14612 387852 14618
rect 387800 14554 387852 14560
rect 387708 5908 387760 5914
rect 387708 5850 387760 5856
rect 386328 5772 386380 5778
rect 386328 5714 386380 5720
rect 387156 4004 387208 4010
rect 387156 3946 387208 3952
rect 387168 480 387196 3946
rect 387812 490 387840 14554
rect 389008 5982 389036 57462
rect 389100 6050 389128 59758
rect 390020 57526 390048 59758
rect 390940 57526 390968 59758
rect 390008 57520 390060 57526
rect 390008 57462 390060 57468
rect 390468 57520 390520 57526
rect 390468 57462 390520 57468
rect 390928 57520 390980 57526
rect 390928 57462 390980 57468
rect 391756 57520 391808 57526
rect 391756 57462 391808 57468
rect 389824 57180 389876 57186
rect 389824 57122 389876 57128
rect 389456 6724 389508 6730
rect 389456 6666 389508 6672
rect 389088 6044 389140 6050
rect 389088 5986 389140 5992
rect 388996 5976 389048 5982
rect 388996 5918 389048 5924
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 6666
rect 389836 5642 389864 57122
rect 390480 6118 390508 57462
rect 391768 6254 391796 57462
rect 391860 6798 391888 59758
rect 392688 57526 392716 59758
rect 393608 57526 393636 59758
rect 392676 57520 392728 57526
rect 392676 57462 392728 57468
rect 393228 57520 393280 57526
rect 393228 57462 393280 57468
rect 393596 57520 393648 57526
rect 393596 57462 393648 57468
rect 394516 57520 394568 57526
rect 394516 57462 394568 57468
rect 391848 6792 391900 6798
rect 391848 6734 391900 6740
rect 393240 6730 393268 57462
rect 393228 6724 393280 6730
rect 393228 6666 393280 6672
rect 394528 6662 394556 57462
rect 393044 6656 393096 6662
rect 393044 6598 393096 6604
rect 394516 6656 394568 6662
rect 394516 6598 394568 6604
rect 391756 6248 391808 6254
rect 391756 6190 391808 6196
rect 390468 6112 390520 6118
rect 390468 6054 390520 6060
rect 389824 5636 389876 5642
rect 389824 5578 389876 5584
rect 391848 5636 391900 5642
rect 391848 5578 391900 5584
rect 390652 4072 390704 4078
rect 390652 4014 390704 4020
rect 390664 480 390692 4014
rect 391860 480 391888 5578
rect 393056 480 393084 6598
rect 394620 6594 394648 59758
rect 395448 57526 395476 59758
rect 396368 57526 396396 59758
rect 395436 57520 395488 57526
rect 395436 57462 395488 57468
rect 395988 57520 396040 57526
rect 395988 57462 396040 57468
rect 396356 57520 396408 57526
rect 396356 57462 396408 57468
rect 394792 57452 394844 57458
rect 394792 57394 394844 57400
rect 394804 54534 394832 57394
rect 394792 54528 394844 54534
rect 394792 54470 394844 54476
rect 394700 24132 394752 24138
rect 394700 24074 394752 24080
rect 394712 16574 394740 24074
rect 394712 16546 395384 16574
rect 394608 6588 394660 6594
rect 394608 6530 394660 6536
rect 394240 4140 394292 4146
rect 394240 4082 394292 4088
rect 394252 480 394280 4082
rect 395356 480 395384 16546
rect 396000 6914 396028 57462
rect 395908 6886 396028 6914
rect 395908 6526 395936 6886
rect 395896 6520 395948 6526
rect 395896 6462 395948 6468
rect 396540 6452 396592 6458
rect 396540 6394 396592 6400
rect 396552 480 396580 6394
rect 397288 6390 397316 59758
rect 398208 57526 398236 59758
rect 399036 57526 399064 59758
rect 397368 57520 397420 57526
rect 397368 57462 397420 57468
rect 398196 57520 398248 57526
rect 398196 57462 398248 57468
rect 398748 57520 398800 57526
rect 398748 57462 398800 57468
rect 399024 57520 399076 57526
rect 399024 57462 399076 57468
rect 397380 6458 397408 57462
rect 397368 6452 397420 6458
rect 397368 6394 397420 6400
rect 397276 6384 397328 6390
rect 397276 6326 397328 6332
rect 398760 6322 398788 57462
rect 398932 13320 398984 13326
rect 398932 13262 398984 13268
rect 398748 6316 398800 6322
rect 398748 6258 398800 6264
rect 397736 3392 397788 3398
rect 397736 3334 397788 3340
rect 397748 480 397776 3334
rect 398944 480 398972 13262
rect 400048 6186 400076 59758
rect 400232 59758 400868 59786
rect 401612 59758 401788 59786
rect 402624 59758 402708 59786
rect 402992 59758 403628 59786
rect 404464 59758 404548 59786
rect 405384 59758 405468 59786
rect 405752 59758 406296 59786
rect 407132 59758 407216 59786
rect 407408 59758 408136 59786
rect 408972 59758 409056 59786
rect 409948 59786 409976 60044
rect 410868 59786 410896 60044
rect 411788 59786 411816 60044
rect 409948 59758 410012 59786
rect 400128 57520 400180 57526
rect 400128 57462 400180 57468
rect 400140 6254 400168 57462
rect 400232 10334 400260 59758
rect 400864 57180 400916 57186
rect 400864 57122 400916 57128
rect 400220 10328 400272 10334
rect 400220 10270 400272 10276
rect 400128 6248 400180 6254
rect 400128 6190 400180 6196
rect 399944 6180 399996 6186
rect 399944 6122 399996 6128
rect 400036 6180 400088 6186
rect 400036 6122 400088 6128
rect 399956 2802 399984 6122
rect 400876 4214 400904 57122
rect 401612 10402 401640 59758
rect 402624 55894 402652 59758
rect 402612 55888 402664 55894
rect 402612 55830 402664 55836
rect 402992 28286 403020 59758
rect 404464 57526 404492 59758
rect 404452 57520 404504 57526
rect 404452 57462 404504 57468
rect 403624 57452 403676 57458
rect 403624 57394 403676 57400
rect 402980 28280 403032 28286
rect 402980 28222 403032 28228
rect 403636 14822 403664 57394
rect 405384 57254 405412 59758
rect 405372 57248 405424 57254
rect 405372 57190 405424 57196
rect 403624 14816 403676 14822
rect 403624 14758 403676 14764
rect 401600 10396 401652 10402
rect 401600 10338 401652 10344
rect 403624 7064 403676 7070
rect 403624 7006 403676 7012
rect 400864 4208 400916 4214
rect 400864 4150 400916 4156
rect 402520 4208 402572 4214
rect 402520 4150 402572 4156
rect 401324 3324 401376 3330
rect 401324 3266 401376 3272
rect 399956 2774 400168 2802
rect 400140 480 400168 2774
rect 401336 480 401364 3266
rect 402532 480 402560 4150
rect 403636 480 403664 7006
rect 405752 3466 405780 59758
rect 407132 57322 407160 59758
rect 407120 57316 407172 57322
rect 407120 57258 407172 57264
rect 405832 31068 405884 31074
rect 405832 31010 405884 31016
rect 405844 16574 405872 31010
rect 407212 18760 407264 18766
rect 407212 18702 407264 18708
rect 405844 16546 406056 16574
rect 405740 3460 405792 3466
rect 405740 3402 405792 3408
rect 404820 3256 404872 3262
rect 404820 3198 404872 3204
rect 404832 480 404860 3198
rect 406028 480 406056 16546
rect 407224 480 407252 18702
rect 407408 3534 407436 59758
rect 408972 57390 409000 59758
rect 408960 57384 409012 57390
rect 408960 57326 409012 57332
rect 409144 11960 409196 11966
rect 409144 11902 409196 11908
rect 407396 3528 407448 3534
rect 407396 3470 407448 3476
rect 408408 3460 408460 3466
rect 408408 3402 408460 3408
rect 408420 480 408448 3402
rect 409156 490 409184 11902
rect 409984 10470 410012 59758
rect 410076 59758 410896 59786
rect 411272 59758 411816 59786
rect 412708 59786 412736 60044
rect 413536 59786 413564 60044
rect 414456 59786 414484 60044
rect 412708 59758 412864 59786
rect 410076 10538 410104 59758
rect 410800 12300 410852 12306
rect 410800 12242 410852 12248
rect 410064 10532 410116 10538
rect 410064 10474 410116 10480
rect 409972 10464 410024 10470
rect 409972 10406 410024 10412
rect 409432 598 409644 626
rect 409432 490 409460 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 462 409460 490
rect 409616 480 409644 598
rect 410812 480 410840 12242
rect 411272 10606 411300 59758
rect 412732 57520 412784 57526
rect 412732 57462 412784 57468
rect 412640 14680 412692 14686
rect 412640 14622 412692 14628
rect 411260 10600 411312 10606
rect 411260 10542 411312 10548
rect 411904 3528 411956 3534
rect 411904 3470 411956 3476
rect 411916 480 411944 3470
rect 412652 490 412680 14622
rect 412744 10742 412772 57462
rect 412732 10736 412784 10742
rect 412732 10678 412784 10684
rect 412836 10674 412864 59758
rect 413480 59758 413564 59786
rect 414032 59758 414484 59786
rect 415376 59786 415404 60044
rect 416296 59786 416324 60044
rect 417216 59786 417244 60044
rect 415376 59758 415532 59786
rect 413480 57526 413508 59758
rect 413468 57520 413520 57526
rect 413468 57462 413520 57468
rect 414032 10810 414060 59758
rect 415400 57520 415452 57526
rect 415400 57462 415452 57468
rect 415412 10946 415440 57462
rect 415400 10940 415452 10946
rect 415400 10882 415452 10888
rect 415504 10878 415532 59758
rect 416240 59758 416324 59786
rect 416792 59758 417244 59786
rect 418136 59786 418164 60044
rect 419056 59786 419084 60044
rect 419976 59786 420004 60044
rect 420804 59786 420832 60044
rect 421724 59786 421752 60044
rect 422644 59786 422672 60044
rect 423564 59786 423592 60044
rect 424484 59786 424512 60044
rect 425404 59786 425432 60044
rect 426324 59786 426352 60044
rect 427244 59786 427272 60044
rect 418136 59758 418292 59786
rect 416240 57526 416268 59758
rect 416228 57520 416280 57526
rect 416228 57462 416280 57468
rect 416688 57248 416740 57254
rect 416688 57190 416740 57196
rect 415492 10872 415544 10878
rect 415492 10814 415544 10820
rect 414020 10804 414072 10810
rect 414020 10746 414072 10752
rect 412824 10668 412876 10674
rect 412824 10610 412876 10616
rect 414296 8424 414348 8430
rect 414296 8366 414348 8372
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 8366
rect 416412 7132 416464 7138
rect 416412 7074 416464 7080
rect 415492 3052 415544 3058
rect 415492 2994 415544 3000
rect 415504 480 415532 2994
rect 416424 2774 416452 7074
rect 416700 3058 416728 57190
rect 416792 11014 416820 59758
rect 418160 57520 418212 57526
rect 418160 57462 418212 57468
rect 416780 11008 416832 11014
rect 416780 10950 416832 10956
rect 418172 10198 418200 57462
rect 418264 10266 418292 59758
rect 419000 59758 419084 59786
rect 419552 59758 420004 59786
rect 420104 59758 420832 59786
rect 420932 59758 421752 59786
rect 422312 59758 422672 59786
rect 422772 59758 423592 59786
rect 423692 59758 424512 59786
rect 425072 59758 425432 59786
rect 425532 59758 426352 59786
rect 427188 59758 427272 59786
rect 427820 59832 427872 59838
rect 428072 59786 428100 60044
rect 428992 59838 429020 60044
rect 427820 59774 427872 59780
rect 419000 57526 419028 59758
rect 418988 57520 419040 57526
rect 418988 57462 419040 57468
rect 418252 10260 418304 10266
rect 418252 10202 418304 10208
rect 418160 10192 418212 10198
rect 418160 10134 418212 10140
rect 419552 10130 419580 59758
rect 420104 45554 420132 59758
rect 419644 45526 420132 45554
rect 419540 10124 419592 10130
rect 419540 10066 419592 10072
rect 419644 10062 419672 45526
rect 419632 10056 419684 10062
rect 419632 9998 419684 10004
rect 420932 9994 420960 59758
rect 421564 57384 421616 57390
rect 421564 57326 421616 57332
rect 421576 18630 421604 57326
rect 421564 18624 421616 18630
rect 421564 18566 421616 18572
rect 420920 9988 420972 9994
rect 420920 9930 420972 9936
rect 422312 9926 422340 59758
rect 422772 45554 422800 59758
rect 423588 57316 423640 57322
rect 423588 57258 423640 57264
rect 422404 45526 422800 45554
rect 422300 9920 422352 9926
rect 422300 9862 422352 9868
rect 422404 9858 422432 45526
rect 422392 9852 422444 9858
rect 422392 9794 422444 9800
rect 421380 8560 421432 8566
rect 421380 8502 421432 8508
rect 417884 8492 417936 8498
rect 417884 8434 417936 8440
rect 416688 3052 416740 3058
rect 416688 2994 416740 3000
rect 416424 2746 416728 2774
rect 416700 480 416728 2746
rect 417896 480 417924 8434
rect 420184 7200 420236 7206
rect 420184 7142 420236 7148
rect 418988 3120 419040 3126
rect 418988 3062 419040 3068
rect 419000 480 419028 3062
rect 420196 480 420224 7142
rect 421392 480 421420 8502
rect 423600 3194 423628 57258
rect 423692 21418 423720 59758
rect 423680 21412 423732 21418
rect 423680 21354 423732 21360
rect 425072 15978 425100 59758
rect 425532 45554 425560 59758
rect 427188 57390 427216 59758
rect 427176 57384 427228 57390
rect 427176 57326 427228 57332
rect 425164 45526 425560 45554
rect 425164 32434 425192 45526
rect 425152 32428 425204 32434
rect 425152 32370 425204 32376
rect 427832 16046 427860 59774
rect 427924 59758 428100 59786
rect 428980 59832 429032 59838
rect 429912 59786 429940 60044
rect 428980 59774 429032 59780
rect 429212 59758 429940 59786
rect 430580 59832 430632 59838
rect 430832 59786 430860 60044
rect 431752 59838 431780 60044
rect 430580 59774 430632 59780
rect 427924 37942 427952 59758
rect 427912 37936 427964 37942
rect 427912 37878 427964 37884
rect 427820 16040 427872 16046
rect 427820 15982 427872 15988
rect 425060 15972 425112 15978
rect 425060 15914 425112 15920
rect 429212 14550 429240 59758
rect 429844 56636 429896 56642
rect 429844 56578 429896 56584
rect 429200 14544 429252 14550
rect 429200 14486 429252 14492
rect 429856 13258 429884 56578
rect 430592 16114 430620 59774
rect 430684 59758 430860 59786
rect 431740 59832 431792 59838
rect 432672 59786 432700 60044
rect 433592 59786 433620 60044
rect 434512 59786 434540 60044
rect 435340 59786 435368 60044
rect 431740 59774 431792 59780
rect 431972 59758 432700 59786
rect 433536 59758 433620 59786
rect 434456 59758 434540 59786
rect 434732 59758 435368 59786
rect 436100 59832 436152 59838
rect 436260 59786 436288 60044
rect 437180 59838 437208 60044
rect 436100 59774 436152 59780
rect 430684 33794 430712 59758
rect 430672 33788 430724 33794
rect 430672 33730 430724 33736
rect 431972 26926 432000 59758
rect 433248 57384 433300 57390
rect 433248 57326 433300 57332
rect 431960 26920 432012 26926
rect 431960 26862 432012 26868
rect 430580 16108 430632 16114
rect 430580 16050 430632 16056
rect 429844 13252 429896 13258
rect 429844 13194 429896 13200
rect 432052 8764 432104 8770
rect 432052 8706 432104 8712
rect 428464 8696 428516 8702
rect 428464 8638 428516 8644
rect 424968 8628 425020 8634
rect 424968 8570 425020 8576
rect 423772 7268 423824 7274
rect 423772 7210 423824 7216
rect 422576 3188 422628 3194
rect 422576 3130 422628 3136
rect 423588 3188 423640 3194
rect 423588 3130 423640 3136
rect 422588 480 422616 3130
rect 423784 480 423812 7210
rect 424980 480 425008 8570
rect 427268 7336 427320 7342
rect 427268 7278 427320 7284
rect 426164 3052 426216 3058
rect 426164 2994 426216 3000
rect 426176 480 426204 2994
rect 427280 480 427308 7278
rect 428476 480 428504 8638
rect 430856 7404 430908 7410
rect 430856 7346 430908 7352
rect 429660 3052 429712 3058
rect 429660 2994 429712 3000
rect 429672 480 429700 2994
rect 430868 480 430896 7346
rect 432064 480 432092 8706
rect 433260 480 433288 57326
rect 433536 56098 433564 59758
rect 434456 56642 434484 59758
rect 434444 56636 434496 56642
rect 434444 56578 434496 56584
rect 433524 56092 433576 56098
rect 433524 56034 433576 56040
rect 434732 17338 434760 59758
rect 435364 57520 435416 57526
rect 435364 57462 435416 57468
rect 434720 17332 434772 17338
rect 434720 17274 434772 17280
rect 435376 13394 435404 57462
rect 436112 17270 436140 59774
rect 436204 59758 436288 59786
rect 437168 59832 437220 59838
rect 438100 59786 438128 60044
rect 437168 59774 437220 59780
rect 438044 59758 438128 59786
rect 438860 59832 438912 59838
rect 439020 59786 439048 60044
rect 439940 59838 439968 60044
rect 438860 59774 438912 59780
rect 436204 25566 436232 59758
rect 438044 57458 438072 59758
rect 438032 57452 438084 57458
rect 438032 57394 438084 57400
rect 436192 25560 436244 25566
rect 436192 25502 436244 25508
rect 436100 17264 436152 17270
rect 436100 17206 436152 17212
rect 438872 14890 438900 59774
rect 438964 59758 439048 59786
rect 439928 59832 439980 59838
rect 440860 59786 440888 60044
rect 441780 59922 441808 60044
rect 439928 59774 439980 59780
rect 440804 59758 440888 59786
rect 441724 59894 441808 59922
rect 438964 29646 438992 59758
rect 440804 57526 440832 59758
rect 440792 57520 440844 57526
rect 440792 57462 440844 57468
rect 441528 57452 441580 57458
rect 441528 57394 441580 57400
rect 438952 29640 439004 29646
rect 438952 29582 439004 29588
rect 438860 14884 438912 14890
rect 438860 14826 438912 14832
rect 435364 13388 435416 13394
rect 435364 13330 435416 13336
rect 439136 8900 439188 8906
rect 439136 8842 439188 8848
rect 435548 8832 435600 8838
rect 435548 8774 435600 8780
rect 434444 7472 434496 7478
rect 434444 7414 434496 7420
rect 434456 480 434484 7414
rect 435560 480 435588 8774
rect 437940 7540 437992 7546
rect 437940 7482 437992 7488
rect 436744 2916 436796 2922
rect 436744 2858 436796 2864
rect 436756 480 436784 2858
rect 437952 480 437980 7482
rect 439148 480 439176 8842
rect 441252 8288 441304 8294
rect 441252 8230 441304 8236
rect 440332 2984 440384 2990
rect 440332 2926 440384 2932
rect 440344 480 440372 2926
rect 441264 2774 441292 8230
rect 441540 2990 441568 57394
rect 441724 56234 441752 59894
rect 442608 59786 442636 60044
rect 443528 59786 443556 60044
rect 444448 59786 444476 60044
rect 445368 59786 445396 60044
rect 446288 59786 446316 60044
rect 441908 59758 442636 59786
rect 443012 59758 443556 59786
rect 444392 59758 444476 59786
rect 445312 59758 445396 59786
rect 445772 59758 446316 59786
rect 447208 59786 447236 60044
rect 448128 59786 448156 60044
rect 449048 59786 449076 60044
rect 447208 59758 447272 59786
rect 441712 56228 441764 56234
rect 441712 56170 441764 56176
rect 441908 45554 441936 59758
rect 441632 45526 441936 45554
rect 441632 35222 441660 45526
rect 441620 35216 441672 35222
rect 441620 35158 441672 35164
rect 443012 19990 443040 59758
rect 443644 57860 443696 57866
rect 443644 57802 443696 57808
rect 443000 19984 443052 19990
rect 443000 19926 443052 19932
rect 442632 9648 442684 9654
rect 442632 9590 442684 9596
rect 441528 2984 441580 2990
rect 441528 2926 441580 2932
rect 441264 2746 441568 2774
rect 441540 480 441568 2746
rect 442644 480 442672 9590
rect 443656 8294 443684 57802
rect 444392 57594 444420 59758
rect 444380 57588 444432 57594
rect 444380 57530 444432 57536
rect 445312 56166 445340 59758
rect 445300 56160 445352 56166
rect 445300 56102 445352 56108
rect 445772 12034 445800 59758
rect 447140 56160 447192 56166
rect 447140 56102 447192 56108
rect 447152 36582 447180 56102
rect 447244 54602 447272 59758
rect 448072 59758 448156 59786
rect 448532 59758 449076 59786
rect 449876 59786 449904 60044
rect 450796 59786 450824 60044
rect 451716 59786 451744 60044
rect 449876 59758 450032 59786
rect 448072 56166 448100 59758
rect 448428 57520 448480 57526
rect 448428 57462 448480 57468
rect 448060 56160 448112 56166
rect 448060 56102 448112 56108
rect 447232 54596 447284 54602
rect 447232 54538 447284 54544
rect 447140 36576 447192 36582
rect 447140 36518 447192 36524
rect 445760 12028 445812 12034
rect 445760 11970 445812 11976
rect 446220 9580 446272 9586
rect 446220 9522 446272 9528
rect 443644 8288 443696 8294
rect 443644 8230 443696 8236
rect 445024 8220 445076 8226
rect 445024 8162 445076 8168
rect 443828 2848 443880 2854
rect 443828 2790 443880 2796
rect 443840 480 443868 2790
rect 445036 480 445064 8162
rect 446232 480 446260 9522
rect 448440 2990 448468 57462
rect 448532 22778 448560 59758
rect 449164 57792 449216 57798
rect 449164 57734 449216 57740
rect 448520 22772 448572 22778
rect 448520 22714 448572 22720
rect 449176 9518 449204 57734
rect 449900 57588 449952 57594
rect 449900 57530 449952 57536
rect 449912 14754 449940 57530
rect 450004 18698 450032 59758
rect 450740 59758 450824 59786
rect 451660 59758 451744 59786
rect 452636 59786 452664 60044
rect 453556 59786 453584 60044
rect 454476 59786 454504 60044
rect 452636 59758 452792 59786
rect 450740 57594 450768 59758
rect 450728 57588 450780 57594
rect 450728 57530 450780 57536
rect 451660 56302 451688 59758
rect 452660 57588 452712 57594
rect 452660 57530 452712 57536
rect 451648 56296 451700 56302
rect 451648 56238 451700 56244
rect 449992 18692 450044 18698
rect 449992 18634 450044 18640
rect 449900 14748 449952 14754
rect 449900 14690 449952 14696
rect 452672 13462 452700 57530
rect 452764 39370 452792 59758
rect 453500 59758 453584 59786
rect 454052 59758 454504 59786
rect 455396 59786 455424 60044
rect 456316 59786 456344 60044
rect 455396 59758 455460 59786
rect 453500 57594 453528 59758
rect 453488 57588 453540 57594
rect 453488 57530 453540 57536
rect 454052 40730 454080 59758
rect 455432 57730 455460 59758
rect 456260 59758 456344 59786
rect 456800 59832 456852 59838
rect 457144 59786 457172 60044
rect 458064 59838 458092 60044
rect 456800 59774 456852 59780
rect 455420 57724 455472 57730
rect 455420 57666 455472 57672
rect 455328 57588 455380 57594
rect 455328 57530 455380 57536
rect 454040 40724 454092 40730
rect 454040 40666 454092 40672
rect 452752 39364 452804 39370
rect 452752 39306 452804 39312
rect 452660 13456 452712 13462
rect 452660 13398 452712 13404
rect 449808 9648 449860 9654
rect 449808 9590 449860 9596
rect 449164 9512 449216 9518
rect 449164 9454 449216 9460
rect 448612 8152 448664 8158
rect 448612 8094 448664 8100
rect 447416 2984 447468 2990
rect 447416 2926 447468 2932
rect 448428 2984 448480 2990
rect 448428 2926 448480 2932
rect 447428 480 447456 2926
rect 448624 480 448652 8094
rect 449820 480 449848 9590
rect 453304 9580 453356 9586
rect 453304 9522 453356 9528
rect 452108 8084 452160 8090
rect 452108 8026 452160 8032
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 450924 480 450952 2790
rect 452120 480 452148 8026
rect 453316 480 453344 9522
rect 455340 3602 455368 57530
rect 456260 56370 456288 59758
rect 456248 56364 456300 56370
rect 456248 56306 456300 56312
rect 455696 8016 455748 8022
rect 455696 7958 455748 7964
rect 454500 3596 454552 3602
rect 454500 3538 454552 3544
rect 455328 3596 455380 3602
rect 455328 3538 455380 3544
rect 454512 480 454540 3538
rect 455708 480 455736 7958
rect 456812 4214 456840 59774
rect 456904 59758 457172 59786
rect 458052 59832 458104 59838
rect 458984 59786 459012 60044
rect 459904 59786 459932 60044
rect 460824 59786 460852 60044
rect 461744 59786 461772 60044
rect 462664 59786 462692 60044
rect 463584 59786 463612 60044
rect 464412 59786 464440 60044
rect 465332 59786 465360 60044
rect 466252 59786 466280 60044
rect 467172 59786 467200 60044
rect 458052 59774 458104 59780
rect 458192 59758 459012 59786
rect 459664 59758 459932 59786
rect 460216 59758 460852 59786
rect 460952 59758 461772 59786
rect 462424 59758 462692 59786
rect 462792 59758 463612 59786
rect 463712 59758 464440 59786
rect 465184 59758 465360 59786
rect 465552 59758 466280 59786
rect 466472 59758 467200 59786
rect 467840 59832 467892 59838
rect 468092 59786 468120 60044
rect 469012 59838 469040 60044
rect 467840 59774 467892 59780
rect 456904 17474 456932 59758
rect 456892 17468 456944 17474
rect 456892 17410 456944 17416
rect 456892 9376 456944 9382
rect 456892 9318 456944 9324
rect 456800 4208 456852 4214
rect 456800 4150 456852 4156
rect 456904 480 456932 9318
rect 458088 3664 458140 3670
rect 458088 3606 458140 3612
rect 458100 480 458128 3606
rect 458192 3369 458220 59758
rect 459192 7948 459244 7954
rect 459192 7890 459244 7896
rect 458178 3360 458234 3369
rect 458178 3295 458234 3304
rect 459204 480 459232 7890
rect 459664 3505 459692 59758
rect 460216 45554 460244 59758
rect 459756 45526 460244 45554
rect 459756 3641 459784 45526
rect 460388 9308 460440 9314
rect 460388 9250 460440 9256
rect 459742 3632 459798 3641
rect 459742 3567 459798 3576
rect 459650 3496 459706 3505
rect 459650 3431 459706 3440
rect 460400 480 460428 9250
rect 460952 3777 460980 59758
rect 462228 57724 462280 57730
rect 462228 57666 462280 57672
rect 460938 3768 460994 3777
rect 460938 3703 460994 3712
rect 460938 3496 460994 3505
rect 462240 3466 462268 57666
rect 462424 3806 462452 59758
rect 462792 45554 462820 59758
rect 462516 45526 462820 45554
rect 462412 3800 462464 3806
rect 462412 3742 462464 3748
rect 462516 3602 462544 45526
rect 462780 7880 462832 7886
rect 462780 7822 462832 7828
rect 462596 3800 462648 3806
rect 462596 3742 462648 3748
rect 462504 3596 462556 3602
rect 462504 3538 462556 3544
rect 462608 3505 462636 3742
rect 462594 3496 462650 3505
rect 460938 3431 460994 3440
rect 461584 3460 461636 3466
rect 460952 3398 460980 3431
rect 461584 3402 461636 3408
rect 462228 3460 462280 3466
rect 462594 3431 462650 3440
rect 462228 3402 462280 3408
rect 460940 3392 460992 3398
rect 460940 3334 460992 3340
rect 461596 480 461624 3402
rect 462792 480 462820 7822
rect 463712 3874 463740 59758
rect 463976 9240 464028 9246
rect 463976 9182 464028 9188
rect 463700 3868 463752 3874
rect 463700 3810 463752 3816
rect 463988 480 464016 9182
rect 465184 4010 465212 59758
rect 465552 45554 465580 59758
rect 466368 57792 466420 57798
rect 466368 57734 466420 57740
rect 465276 45526 465580 45554
rect 465172 4004 465224 4010
rect 465172 3946 465224 3952
rect 465276 3942 465304 45526
rect 466276 7812 466328 7818
rect 466276 7754 466328 7760
rect 465264 3936 465316 3942
rect 465264 3878 465316 3884
rect 465172 3460 465224 3466
rect 465172 3402 465224 3408
rect 465184 480 465212 3402
rect 466288 480 466316 7754
rect 466380 3466 466408 57734
rect 466472 4078 466500 59758
rect 467104 13592 467156 13598
rect 467104 13534 467156 13540
rect 466460 4072 466512 4078
rect 466460 4014 466512 4020
rect 467116 3602 467144 13534
rect 467472 9172 467524 9178
rect 467472 9114 467524 9120
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 466368 3460 466420 3466
rect 466368 3402 466420 3408
rect 467484 480 467512 9114
rect 467852 4146 467880 59774
rect 467944 59758 468120 59786
rect 469000 59832 469052 59838
rect 469932 59786 469960 60044
rect 470852 59786 470880 60044
rect 471680 59786 471708 60044
rect 472600 59786 472628 60044
rect 469000 59774 469052 59780
rect 469232 59758 469960 59786
rect 470704 59758 470880 59786
rect 470980 59758 471708 59786
rect 472084 59758 472628 59786
rect 473520 59786 473548 60044
rect 474440 59786 474468 60044
rect 475360 59786 475388 60044
rect 476280 59922 476308 60044
rect 473520 59758 473584 59786
rect 467840 4140 467892 4146
rect 467840 4082 467892 4088
rect 467944 3398 467972 59758
rect 469128 57928 469180 57934
rect 469128 57870 469180 57876
rect 469140 3466 469168 57870
rect 469232 3806 469260 59758
rect 469864 7744 469916 7750
rect 469864 7686 469916 7692
rect 469220 3800 469272 3806
rect 469220 3742 469272 3748
rect 468668 3460 468720 3466
rect 468668 3402 468720 3408
rect 469128 3460 469180 3466
rect 469128 3402 469180 3408
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 468680 480 468708 3402
rect 469876 480 469904 7686
rect 470704 3330 470732 59758
rect 470980 45554 471008 59758
rect 470796 45526 471008 45554
rect 470692 3324 470744 3330
rect 470692 3266 470744 3272
rect 470796 3262 470824 45526
rect 471060 9104 471112 9110
rect 471060 9046 471112 9052
rect 470784 3256 470836 3262
rect 470784 3198 470836 3204
rect 471072 480 471100 9046
rect 472084 3738 472112 59758
rect 473268 57860 473320 57866
rect 473268 57802 473320 57808
rect 472072 3732 472124 3738
rect 472072 3674 472124 3680
rect 473280 3534 473308 57802
rect 473452 7676 473504 7682
rect 473452 7618 473504 7624
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 473268 3528 473320 3534
rect 473268 3470 473320 3476
rect 472268 480 472296 3470
rect 473464 480 473492 7618
rect 473556 3466 473584 59758
rect 474384 59758 474468 59786
rect 474844 59758 475388 59786
rect 476224 59894 476308 59922
rect 474384 57254 474412 59758
rect 474372 57248 474424 57254
rect 474372 57190 474424 57196
rect 474556 9036 474608 9042
rect 474556 8978 474608 8984
rect 473544 3460 473596 3466
rect 473544 3402 473596 3408
rect 474568 480 474596 8978
rect 474844 3194 474872 59758
rect 476224 57322 476252 59894
rect 477200 59786 477228 60044
rect 478120 59786 478148 60044
rect 478948 59922 478976 60044
rect 476316 59758 477228 59786
rect 477512 59758 478148 59786
rect 478892 59894 478976 59922
rect 476212 57316 476264 57322
rect 476212 57258 476264 57264
rect 476028 57248 476080 57254
rect 476028 57190 476080 57196
rect 476040 6914 476068 57190
rect 475764 6886 476068 6914
rect 474832 3188 474884 3194
rect 474832 3130 474884 3136
rect 475764 480 475792 6886
rect 476316 3126 476344 59758
rect 476948 7608 477000 7614
rect 476948 7550 477000 7556
rect 476304 3120 476356 3126
rect 476304 3062 476356 3068
rect 476960 480 476988 7550
rect 477512 3058 477540 59758
rect 478892 57390 478920 59894
rect 479868 59786 479896 60044
rect 480788 59786 480816 60044
rect 478984 59758 479896 59786
rect 480732 59758 480816 59786
rect 481708 59786 481736 60044
rect 482628 59786 482656 60044
rect 483548 59786 483576 60044
rect 484468 59786 484496 60044
rect 485388 59786 485416 60044
rect 486308 59786 486336 60044
rect 481708 59758 481864 59786
rect 478880 57384 478932 57390
rect 478880 57326 478932 57332
rect 478144 8968 478196 8974
rect 478144 8910 478196 8916
rect 477500 3052 477552 3058
rect 477500 2994 477552 3000
rect 478156 480 478184 8910
rect 478984 2990 479012 59758
rect 480732 57458 480760 59758
rect 480720 57452 480772 57458
rect 480720 57394 480772 57400
rect 480168 57384 480220 57390
rect 480168 57326 480220 57332
rect 480180 3534 480208 57326
rect 480536 11892 480588 11898
rect 480536 11834 480588 11840
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 478972 2984 479024 2990
rect 478972 2926 479024 2932
rect 479352 480 479380 3470
rect 480548 480 480576 11834
rect 481732 8288 481784 8294
rect 481732 8230 481784 8236
rect 481744 480 481772 8230
rect 481836 2922 481864 59758
rect 482572 59758 482656 59786
rect 483032 59758 483576 59786
rect 484412 59758 484496 59786
rect 484596 59758 485416 59786
rect 486252 59758 486336 59786
rect 487136 59786 487164 60044
rect 488056 59786 488084 60044
rect 488976 59786 489004 60044
rect 487136 59758 487200 59786
rect 482572 57526 482600 59758
rect 482560 57520 482612 57526
rect 482560 57462 482612 57468
rect 482928 57316 482980 57322
rect 482928 57258 482980 57264
rect 482940 6914 482968 57258
rect 482848 6886 482968 6914
rect 481824 2916 481876 2922
rect 481824 2858 481876 2864
rect 482848 480 482876 6886
rect 483032 2854 483060 59758
rect 483664 57656 483716 57662
rect 483664 57598 483716 57604
rect 483676 16574 483704 57598
rect 484412 57594 484440 59758
rect 484400 57588 484452 57594
rect 484400 57530 484452 57536
rect 483676 16546 483796 16574
rect 483664 11756 483716 11762
rect 483664 11698 483716 11704
rect 483676 3482 483704 11698
rect 483768 3738 483796 16546
rect 484492 12232 484544 12238
rect 484492 12174 484544 12180
rect 483756 3732 483808 3738
rect 483756 3674 483808 3680
rect 483676 3454 484072 3482
rect 483020 2848 483072 2854
rect 483020 2790 483072 2796
rect 484044 480 484072 3454
rect 484504 1714 484532 12174
rect 484596 3670 484624 59758
rect 486252 57730 486280 59758
rect 487172 57798 487200 59758
rect 488000 59758 488084 59786
rect 488920 59758 489004 59786
rect 489896 59786 489924 60044
rect 490816 59786 490844 60044
rect 491736 59786 491764 60044
rect 489896 59758 489960 59786
rect 488000 57934 488028 59758
rect 487988 57928 488040 57934
rect 487988 57870 488040 57876
rect 488920 57866 488948 59758
rect 488908 57860 488960 57866
rect 488908 57802 488960 57808
rect 487160 57792 487212 57798
rect 487160 57734 487212 57740
rect 486240 57724 486292 57730
rect 486240 57666 486292 57672
rect 487068 57452 487120 57458
rect 487068 57394 487120 57400
rect 486424 17400 486476 17406
rect 486424 17342 486476 17348
rect 486436 16574 486464 17342
rect 486436 16546 486556 16574
rect 484584 3664 484636 3670
rect 484584 3606 484636 3612
rect 486424 3528 486476 3534
rect 486424 3470 486476 3476
rect 484504 1686 484808 1714
rect 484780 490 484808 1686
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 3470
rect 486528 3466 486556 16546
rect 487080 3534 487108 57394
rect 489932 57254 489960 59758
rect 490760 59758 490844 59786
rect 491680 59758 491764 59786
rect 492656 59786 492684 60044
rect 493576 59786 493604 60044
rect 494404 59786 494432 60044
rect 492656 59758 492720 59786
rect 490760 57390 490788 59758
rect 491680 57390 491708 59758
rect 492692 57458 492720 59758
rect 493520 59758 493604 59786
rect 494072 59758 494432 59786
rect 495324 59786 495352 60044
rect 496244 59786 496272 60044
rect 497164 59786 497192 60044
rect 498084 59786 498112 60044
rect 495324 59758 495388 59786
rect 496244 59758 496308 59786
rect 497164 59758 497228 59786
rect 492680 57452 492732 57458
rect 492680 57394 492732 57400
rect 490748 57384 490800 57390
rect 490748 57326 490800 57332
rect 491668 57384 491720 57390
rect 491668 57326 491720 57332
rect 493520 57322 493548 59758
rect 494072 57644 494100 59758
rect 493980 57616 494100 57644
rect 491208 57316 491260 57322
rect 491208 57258 491260 57264
rect 493508 57316 493560 57322
rect 493508 57258 493560 57264
rect 489920 57248 489972 57254
rect 489920 57190 489972 57196
rect 489184 56024 489236 56030
rect 489184 55966 489236 55972
rect 488816 13524 488868 13530
rect 488816 13466 488868 13472
rect 487160 11824 487212 11830
rect 487160 11766 487212 11772
rect 487068 3528 487120 3534
rect 487068 3470 487120 3476
rect 486516 3460 486568 3466
rect 486516 3402 486568 3408
rect 487172 490 487200 11766
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 13466
rect 489196 4078 489224 55966
rect 490564 14476 490616 14482
rect 490564 14418 490616 14424
rect 489184 4072 489236 4078
rect 489184 4014 489236 4020
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 489932 480 489960 3334
rect 490576 3058 490604 14418
rect 491116 4072 491168 4078
rect 491116 4014 491168 4020
rect 490564 3052 490616 3058
rect 490564 2994 490616 3000
rect 491128 480 491156 4014
rect 491220 3398 491248 57258
rect 493324 13116 493376 13122
rect 493324 13058 493376 13064
rect 493336 3466 493364 13058
rect 493980 3534 494008 57616
rect 493508 3528 493560 3534
rect 493508 3470 493560 3476
rect 493968 3528 494020 3534
rect 493968 3470 494020 3476
rect 492312 3460 492364 3466
rect 492312 3402 492364 3408
rect 493324 3460 493376 3466
rect 493324 3402 493376 3408
rect 491208 3392 491260 3398
rect 491208 3334 491260 3340
rect 492324 480 492352 3402
rect 493520 480 493548 3470
rect 494704 3460 494756 3466
rect 494704 3402 494756 3408
rect 494716 480 494744 3402
rect 495360 3330 495388 59758
rect 496280 57662 496308 59758
rect 496268 57656 496320 57662
rect 496268 57598 496320 57604
rect 497200 57594 497228 59758
rect 498028 59758 498112 59786
rect 499004 59786 499032 60044
rect 499924 59786 499952 60044
rect 500844 59786 500872 60044
rect 501672 59786 501700 60044
rect 502592 59786 502620 60044
rect 503512 59786 503540 60044
rect 504432 59786 504460 60044
rect 505352 59786 505380 60044
rect 506272 59786 506300 60044
rect 507192 59786 507220 60044
rect 508112 59786 508140 60044
rect 508940 59786 508968 60044
rect 509860 59786 509888 60044
rect 510780 59786 510808 60044
rect 511700 59786 511728 60044
rect 512620 59786 512648 60044
rect 513540 59786 513568 60044
rect 514460 59786 514488 60044
rect 515380 59786 515408 60044
rect 516208 59786 516236 60044
rect 499004 59758 499068 59786
rect 499924 59758 499988 59786
rect 500844 59758 500908 59786
rect 501672 59758 501736 59786
rect 502592 59758 502656 59786
rect 503512 59758 503576 59786
rect 504432 59758 504496 59786
rect 505352 59758 505416 59786
rect 506272 59758 506336 59786
rect 507192 59758 507256 59786
rect 508112 59758 508176 59786
rect 508940 59758 509188 59786
rect 509860 59758 509924 59786
rect 510780 59758 510844 59786
rect 511700 59758 511948 59786
rect 512620 59758 512684 59786
rect 513540 59758 513604 59786
rect 514460 59758 514616 59786
rect 515380 59758 515444 59786
rect 516208 59758 516272 59786
rect 497464 57656 497516 57662
rect 497464 57598 497516 57604
rect 497188 57588 497240 57594
rect 497188 57530 497240 57536
rect 495440 12164 495492 12170
rect 495440 12106 495492 12112
rect 495348 3324 495400 3330
rect 495348 3266 495400 3272
rect 495452 490 495480 12106
rect 497476 4010 497504 57598
rect 497464 4004 497516 4010
rect 497464 3946 497516 3952
rect 498028 3670 498056 59758
rect 499040 57662 499068 59758
rect 499960 57662 499988 59758
rect 499028 57656 499080 57662
rect 499028 57598 499080 57604
rect 499488 57656 499540 57662
rect 499488 57598 499540 57604
rect 499948 57656 500000 57662
rect 499948 57598 500000 57604
rect 500776 57656 500828 57662
rect 500776 57598 500828 57604
rect 498108 57588 498160 57594
rect 498108 57530 498160 57536
rect 498120 3806 498148 57530
rect 498108 3800 498160 3806
rect 498108 3742 498160 3748
rect 498016 3664 498068 3670
rect 498016 3606 498068 3612
rect 499500 3398 499528 57598
rect 500592 4004 500644 4010
rect 500592 3946 500644 3952
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499488 3392 499540 3398
rect 499488 3334 499540 3340
rect 497096 3324 497148 3330
rect 497096 3266 497148 3272
rect 495728 598 495940 626
rect 495728 490 495756 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 462 495756 490
rect 495912 480 495940 598
rect 497108 480 497136 3266
rect 498200 3052 498252 3058
rect 498200 2994 498252 3000
rect 498212 480 498240 2994
rect 499408 480 499436 3334
rect 500604 480 500632 3946
rect 500788 3466 500816 57598
rect 500776 3460 500828 3466
rect 500776 3402 500828 3408
rect 500880 2990 500908 59758
rect 501708 57458 501736 59758
rect 502628 57662 502656 59758
rect 502616 57656 502668 57662
rect 502616 57598 502668 57604
rect 501696 57452 501748 57458
rect 501696 57394 501748 57400
rect 502248 57452 502300 57458
rect 502248 57394 502300 57400
rect 501328 13184 501380 13190
rect 501328 13126 501380 13132
rect 500868 2984 500920 2990
rect 500868 2926 500920 2932
rect 501340 490 501368 13126
rect 502260 3058 502288 57394
rect 502984 9512 503036 9518
rect 502984 9454 503036 9460
rect 502248 3052 502300 3058
rect 502248 2994 502300 3000
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 9454
rect 503548 3738 503576 59758
rect 503628 57656 503680 57662
rect 503628 57598 503680 57604
rect 503536 3732 503588 3738
rect 503536 3674 503588 3680
rect 503640 3126 503668 57598
rect 504468 57458 504496 59758
rect 505388 57662 505416 59758
rect 505376 57656 505428 57662
rect 505376 57598 505428 57604
rect 504456 57452 504508 57458
rect 504456 57394 504508 57400
rect 505008 57452 505060 57458
rect 505008 57394 505060 57400
rect 504364 55956 504416 55962
rect 504364 55898 504416 55904
rect 504180 3800 504232 3806
rect 504180 3742 504232 3748
rect 503628 3120 503680 3126
rect 503628 3062 503680 3068
rect 504192 480 504220 3742
rect 504376 3534 504404 55898
rect 504364 3528 504416 3534
rect 504364 3470 504416 3476
rect 505020 3194 505048 57394
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 505008 3188 505060 3194
rect 505008 3130 505060 3136
rect 505388 480 505416 3470
rect 506308 3262 506336 59758
rect 506388 57656 506440 57662
rect 506388 57598 506440 57604
rect 506400 3330 506428 57598
rect 507228 57458 507256 59758
rect 508148 57662 508176 59758
rect 508136 57656 508188 57662
rect 508136 57598 508188 57604
rect 509056 57656 509108 57662
rect 509056 57598 509108 57604
rect 507216 57452 507268 57458
rect 507216 57394 507268 57400
rect 507768 57452 507820 57458
rect 507768 57394 507820 57400
rect 507124 15904 507176 15910
rect 507124 15846 507176 15852
rect 506480 12096 506532 12102
rect 506480 12038 506532 12044
rect 506388 3324 506440 3330
rect 506388 3266 506440 3272
rect 506296 3256 506348 3262
rect 506296 3198 506348 3204
rect 506492 480 506520 12038
rect 507136 3534 507164 15846
rect 507780 4146 507808 57394
rect 507768 4140 507820 4146
rect 507768 4082 507820 4088
rect 509068 4078 509096 57598
rect 509056 4072 509108 4078
rect 509056 4014 509108 4020
rect 509160 4010 509188 59758
rect 509896 57662 509924 59758
rect 510816 57662 510844 59758
rect 509884 57656 509936 57662
rect 509884 57598 509936 57604
rect 510528 57656 510580 57662
rect 510528 57598 510580 57604
rect 510804 57656 510856 57662
rect 510804 57598 510856 57604
rect 511816 57656 511868 57662
rect 511816 57598 511868 57604
rect 509148 4004 509200 4010
rect 509148 3946 509200 3952
rect 507676 3664 507728 3670
rect 507676 3606 507728 3612
rect 507124 3528 507176 3534
rect 507124 3470 507176 3476
rect 507688 480 507716 3606
rect 510540 3602 510568 57598
rect 511828 3874 511856 57598
rect 511920 3942 511948 59758
rect 512656 57662 512684 59758
rect 513576 57662 513604 59758
rect 512644 57656 512696 57662
rect 512644 57598 512696 57604
rect 513288 57656 513340 57662
rect 513288 57598 513340 57604
rect 513564 57656 513616 57662
rect 513564 57598 513616 57604
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 511908 3936 511960 3942
rect 511908 3878 511960 3884
rect 511816 3868 511868 3874
rect 511816 3810 511868 3816
rect 510068 3596 510120 3602
rect 510068 3538 510120 3544
rect 510528 3596 510580 3602
rect 510528 3538 510580 3544
rect 508872 3528 508924 3534
rect 508872 3470 508924 3476
rect 508884 480 508912 3470
rect 510080 480 510108 3538
rect 511264 3392 511316 3398
rect 511264 3334 511316 3340
rect 511276 480 511304 3334
rect 512472 480 512500 4218
rect 513300 3806 513328 57598
rect 513564 5636 513616 5642
rect 513564 5578 513616 5584
rect 513288 3800 513340 3806
rect 513288 3742 513340 3748
rect 513576 480 513604 5578
rect 514588 3534 514616 59758
rect 515416 57662 515444 59758
rect 514668 57656 514720 57662
rect 514668 57598 514720 57604
rect 515404 57656 515456 57662
rect 515404 57598 515456 57604
rect 516048 57656 516100 57662
rect 516048 57598 516100 57604
rect 514680 3670 514708 57598
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 514668 3664 514720 3670
rect 514668 3606 514720 3612
rect 514576 3528 514628 3534
rect 514576 3470 514628 3476
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 4286
rect 516060 3534 516088 57598
rect 516244 57594 516272 59758
rect 516232 57588 516284 57594
rect 516232 57530 516284 57536
rect 517428 57588 517480 57594
rect 517428 57530 517480 57536
rect 517152 5704 517204 5710
rect 517152 5646 517204 5652
rect 516048 3528 516100 3534
rect 516048 3470 516100 3476
rect 517164 480 517192 5646
rect 517440 3466 517468 57530
rect 522316 6866 522344 60823
rect 522408 20670 522436 71295
rect 522500 33114 522528 82719
rect 522592 46918 522620 94007
rect 522684 60722 522712 105431
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 522672 60716 522724 60722
rect 522672 60658 522724 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 522580 46912 522632 46918
rect 522580 46854 522632 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 522488 33108 522540 33114
rect 580170 33079 580172 33088
rect 522488 33050 522540 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 522396 20664 522448 20670
rect 522396 20606 522448 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 522304 6860 522356 6866
rect 522304 6802 522356 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 545488 6792 545540 6798
rect 545488 6734 545540 6740
rect 538404 6112 538456 6118
rect 538404 6054 538456 6060
rect 534908 6044 534960 6050
rect 534908 5986 534960 5992
rect 531320 5976 531372 5982
rect 531320 5918 531372 5924
rect 527824 5908 527876 5914
rect 527824 5850 527876 5856
rect 524236 5840 524288 5846
rect 524236 5782 524288 5788
rect 520740 5772 520792 5778
rect 520740 5714 520792 5720
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 517428 3460 517480 3466
rect 517428 3402 517480 3408
rect 518348 2984 518400 2990
rect 518348 2926 518400 2932
rect 518360 480 518388 2926
rect 519556 480 519584 4354
rect 520752 480 520780 5714
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 521844 3052 521896 3058
rect 521844 2994 521896 3000
rect 521856 480 521884 2994
rect 523052 480 523080 4422
rect 524248 480 524276 5782
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 525432 3120 525484 3126
rect 525432 3062 525484 3068
rect 525444 480 525472 3062
rect 526640 480 526668 4490
rect 527836 480 527864 5850
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 529020 3188 529072 3194
rect 529020 3130 529072 3136
rect 529032 480 529060 3130
rect 530136 480 530164 4558
rect 531332 480 531360 5918
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 3256 532568 3262
rect 532516 3198 532568 3204
rect 532528 480 532556 3198
rect 533724 480 533752 4626
rect 534920 480 534948 5986
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 536104 3324 536156 3330
rect 536104 3266 536156 3272
rect 536116 480 536144 3266
rect 537220 480 537248 4694
rect 538416 480 538444 6054
rect 541992 5568 542044 5574
rect 541992 5510 542044 5516
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3392 539652 3398
rect 539600 3334 539652 3340
rect 539612 480 539640 3334
rect 540808 480 540836 5442
rect 542004 480 542032 5510
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 4140 543240 4146
rect 543188 4082 543240 4088
rect 543200 480 543228 4082
rect 544396 480 544424 5374
rect 545500 480 545528 6734
rect 549076 6724 549128 6730
rect 549076 6666 549128 6672
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 4072 546736 4078
rect 546684 4014 546736 4020
rect 546696 480 546724 4014
rect 547892 480 547920 5306
rect 549088 480 549116 6666
rect 552664 6656 552716 6662
rect 580184 6633 580212 6802
rect 552664 6598 552716 6604
rect 580170 6624 580226 6633
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 4004 550324 4010
rect 550272 3946 550324 3952
rect 550284 480 550312 3946
rect 551480 480 551508 5238
rect 552676 480 552704 6598
rect 556160 6588 556212 6594
rect 580170 6559 580226 6568
rect 556160 6530 556212 6536
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3936 553820 3942
rect 553768 3878 553820 3884
rect 553780 480 553808 3878
rect 554976 480 555004 5170
rect 556172 480 556200 6530
rect 559748 6520 559800 6526
rect 559748 6462 559800 6468
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3868 557408 3874
rect 557356 3810 557408 3816
rect 557368 480 557396 3810
rect 558564 480 558592 5102
rect 559760 480 559788 6462
rect 563244 6452 563296 6458
rect 563244 6394 563296 6400
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560852 3800 560904 3806
rect 560852 3742 560904 3748
rect 560864 480 560892 3742
rect 562060 480 562088 5034
rect 563256 480 563284 6394
rect 566832 6384 566884 6390
rect 566832 6326 566884 6332
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3732 564492 3738
rect 564440 3674 564492 3680
rect 564452 480 564480 3674
rect 565648 480 565676 4966
rect 566844 480 566872 6326
rect 570328 6316 570380 6322
rect 570328 6258 570380 6264
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4898
rect 570340 480 570368 6258
rect 573916 6248 573968 6254
rect 573916 6190 573968 6196
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 571536 480 571564 3538
rect 572732 480 572760 4830
rect 573928 480 573956 6190
rect 577412 6180 577464 6186
rect 577412 6122 577464 6128
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3528 575164 3534
rect 575112 3470 575164 3476
rect 575124 480 575152 3470
rect 576320 480 576348 4762
rect 577424 480 577452 6122
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 632032 3478 632088
rect 3606 658144 3662 658200
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 522302 650800 522358 650856
rect 69018 640872 69074 640928
rect 69018 629720 69074 629776
rect 3514 619112 3570 619168
rect 69018 618568 69074 618624
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 522394 640464 522450 640520
rect 522302 606464 522358 606520
rect 3606 606056 3662 606112
rect 3422 579944 3478 580000
rect 69018 596264 69074 596320
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 522486 629176 522542 629232
rect 580170 617480 580226 617536
rect 522394 595040 522450 595096
rect 69018 584976 69074 585032
rect 69018 573824 69074 573880
rect 3514 566888 3570 566944
rect 579802 590960 579858 591016
rect 522486 583616 522542 583672
rect 580170 577632 580226 577688
rect 522302 560768 522358 560824
rect 3606 553832 3662 553888
rect 69018 551520 69074 551576
rect 579802 564304 579858 564360
rect 522394 549480 522450 549536
rect 69018 540368 69074 540424
rect 522486 538056 522542 538112
rect 580170 537784 580226 537840
rect 69018 529216 69074 529272
rect 3422 527856 3478 527912
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 522302 515344 522358 515400
rect 3514 514800 3570 514856
rect 3422 501744 3478 501800
rect 69018 506912 69074 506968
rect 69018 495624 69074 495680
rect 580170 511264 580226 511320
rect 522394 503920 522450 503976
rect 522302 492496 522358 492552
rect 580170 484608 580226 484664
rect 69018 484472 69074 484528
rect 3422 475632 3478 475688
rect 579986 471416 580042 471472
rect 522302 469784 522358 469840
rect 3514 462576 3570 462632
rect 69018 462168 69074 462224
rect 522394 458360 522450 458416
rect 580170 458088 580226 458144
rect 69018 451016 69074 451072
rect 3422 449520 3478 449576
rect 522302 446936 522358 446992
rect 69018 439864 69074 439920
rect 580170 431568 580226 431624
rect 522946 424224 523002 424280
rect 3330 423544 3386 423600
rect 580170 418240 580226 418296
rect 69018 417424 69074 417480
rect 522946 412800 523002 412856
rect 3422 410488 3478 410544
rect 69018 406408 69074 406464
rect 580170 404912 580226 404968
rect 522026 401512 522082 401568
rect 2870 397432 2926 397488
rect 69018 395120 69074 395176
rect 522946 378664 523002 378720
rect 580170 378392 580226 378448
rect 69018 372816 69074 372872
rect 3422 371320 3478 371376
rect 522946 367240 523002 367296
rect 580170 365064 580226 365120
rect 69018 361664 69074 361720
rect 3422 358400 3478 358456
rect 522946 355952 523002 356008
rect 580170 351872 580226 351928
rect 69018 350376 69074 350432
rect 2870 345344 2926 345400
rect 522302 333104 522358 333160
rect 69018 328072 69074 328128
rect 580170 325216 580226 325272
rect 522302 321816 522358 321872
rect 2870 319232 2926 319288
rect 69018 316920 69074 316976
rect 580170 312024 580226 312080
rect 522302 310256 522358 310312
rect 3514 306176 3570 306232
rect 69018 305768 69074 305824
rect 580170 298696 580226 298752
rect 3422 293120 3478 293176
rect 522394 287680 522450 287736
rect 69018 283328 69074 283384
rect 522302 276120 522358 276176
rect 69018 272312 69074 272368
rect 3422 267144 3478 267200
rect 69018 261024 69074 261080
rect 580170 272176 580226 272232
rect 522394 264832 522450 264888
rect 3514 254088 3570 254144
rect 522302 253408 522358 253464
rect 3422 241032 3478 241088
rect 69018 238756 69020 238776
rect 69020 238756 69072 238776
rect 69072 238756 69074 238776
rect 69018 238720 69074 238756
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 522394 241984 522450 242040
rect 522302 230696 522358 230752
rect 69018 227568 69074 227624
rect 3514 214920 3570 214976
rect 69018 216416 69074 216472
rect 579986 232328 580042 232384
rect 522486 219272 522542 219328
rect 522394 207848 522450 207904
rect 3606 201864 3662 201920
rect 522302 196424 522358 196480
rect 69018 194112 69074 194168
rect 3422 188808 3478 188864
rect 69018 182824 69074 182880
rect 69018 171672 69074 171728
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 522486 185136 522542 185192
rect 522394 173848 522450 173904
rect 3606 162832 3662 162888
rect 522302 162288 522358 162344
rect 3514 149776 3570 149832
rect 69018 149368 69074 149424
rect 3422 136720 3478 136776
rect 69018 138216 69074 138272
rect 69018 127064 69074 127120
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 522578 151000 522634 151056
rect 522486 139576 522542 139632
rect 522394 128152 522450 128208
rect 522302 116864 522358 116920
rect 69018 115776 69074 115832
rect 3698 110608 3754 110664
rect 69018 104760 69074 104816
rect 3606 97552 3662 97608
rect 3514 84632 3570 84688
rect 3422 71576 3478 71632
rect 69018 93472 69074 93528
rect 69018 82320 69074 82376
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 522670 105440 522726 105496
rect 522578 94016 522634 94072
rect 522486 82728 522542 82784
rect 522394 71304 522450 71360
rect 69018 71168 69074 71224
rect 69018 61104 69074 61160
rect 522302 60832 522358 60888
rect 3790 58520 3846 58576
rect 3698 45464 3754 45520
rect 3606 32408 3662 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 355230 3304 355286 3360
rect 358726 3440 358782 3496
rect 362314 3576 362370 3632
rect 365810 3712 365866 3768
rect 458178 3304 458234 3360
rect 459742 3576 459798 3632
rect 459650 3440 459706 3496
rect 460938 3712 460994 3768
rect 460938 3440 460994 3496
rect 462594 3440 462650 3496
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3601 658202 3667 658205
rect -960 658200 3667 658202
rect -960 658144 3606 658200
rect 3662 658144 3667 658200
rect -960 658142 3667 658144
rect -960 658052 480 658142
rect 3601 658139 3667 658142
rect 583520 657236 584960 657476
rect 519892 650858 520474 650896
rect 522297 650858 522363 650861
rect 519892 650856 522363 650858
rect 519892 650836 522302 650856
rect 520414 650800 522302 650836
rect 522358 650800 522363 650856
rect 520414 650798 522363 650800
rect 522297 650795 522363 650798
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 69013 640930 69079 640933
rect 69013 640928 71514 640930
rect 69013 640872 69018 640928
rect 69074 640892 71514 640928
rect 69074 640872 72036 640892
rect 69013 640870 72036 640872
rect 69013 640867 69079 640870
rect 71454 640832 72036 640870
rect 519892 640522 520474 640526
rect 522389 640522 522455 640525
rect 519892 640520 522455 640522
rect 519892 640466 522394 640520
rect 520414 640464 522394 640466
rect 522450 640464 522455 640520
rect 520414 640462 522455 640464
rect 522389 640459 522455 640462
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 69013 629778 69079 629781
rect 71454 629778 72036 629790
rect 69013 629776 72036 629778
rect 69013 629720 69018 629776
rect 69074 629730 72036 629776
rect 69074 629720 71514 629730
rect 69013 629718 71514 629720
rect 69013 629715 69079 629718
rect 522481 629234 522547 629237
rect 520414 629232 522547 629234
rect 520414 629180 522486 629232
rect 519892 629176 522486 629180
rect 522542 629176 522547 629232
rect 519892 629174 522547 629176
rect 519892 629120 520474 629174
rect 522481 629171 522547 629174
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 69013 618626 69079 618629
rect 69013 618624 71514 618626
rect 69013 618568 69018 618624
rect 69074 618568 71514 618624
rect 69013 618566 71514 618568
rect 69013 618563 69079 618566
rect 71454 618506 72036 618566
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 522297 606522 522363 606525
rect 520414 606520 522363 606522
rect 520414 606488 522302 606520
rect 519892 606464 522302 606488
rect 522358 606464 522363 606520
rect 519892 606462 522363 606464
rect 519892 606428 520474 606462
rect 522297 606459 522363 606462
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect 69013 596322 69079 596325
rect 69013 596320 71514 596322
rect 69013 596264 69018 596320
rect 69074 596264 71514 596320
rect 69013 596262 71514 596264
rect 69013 596259 69079 596262
rect 71454 596240 71514 596262
rect 71454 596180 72036 596240
rect 522389 595098 522455 595101
rect 520414 595096 522455 595098
rect 520414 595040 522394 595096
rect 522450 595040 522455 595096
rect 520414 595038 522455 595040
rect 520414 595020 520474 595038
rect 522389 595035 522455 595038
rect 519892 594960 520474 595020
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 69013 585034 69079 585037
rect 69013 585032 71514 585034
rect 69013 584976 69018 585032
rect 69074 585016 71514 585032
rect 69074 584976 72036 585016
rect 69013 584974 72036 584976
rect 69013 584971 69079 584974
rect 71454 584956 72036 584974
rect 522481 583674 522547 583677
rect 519892 583672 522547 583674
rect 519892 583616 522486 583672
rect 522542 583616 522547 583672
rect 519892 583614 522547 583616
rect 522481 583611 522547 583614
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 69013 573882 69079 573885
rect 71454 573882 72036 573914
rect 69013 573880 72036 573882
rect 69013 573824 69018 573880
rect 69074 573854 72036 573880
rect 69074 573824 71514 573854
rect 69013 573822 71514 573824
rect 69013 573819 69079 573822
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 519892 560826 520474 560860
rect 522297 560826 522363 560829
rect 519892 560824 522363 560826
rect 519892 560800 522302 560824
rect 520414 560768 522302 560800
rect 522358 560768 522363 560824
rect 520414 560766 522363 560768
rect 522297 560763 522363 560766
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 69013 551578 69079 551581
rect 71454 551578 72036 551588
rect 69013 551576 72036 551578
rect 69013 551520 69018 551576
rect 69074 551528 72036 551576
rect 69074 551520 71514 551528
rect 69013 551518 71514 551520
rect 69013 551515 69079 551518
rect 583520 551020 584960 551260
rect 522389 549538 522455 549541
rect 520414 549536 522455 549538
rect 520414 549514 522394 549536
rect 519892 549480 522394 549514
rect 522450 549480 522455 549536
rect 519892 549478 522455 549480
rect 519892 549454 520474 549478
rect 522389 549475 522455 549478
rect -960 540684 480 540924
rect 69013 540426 69079 540429
rect 69013 540424 71514 540426
rect 69013 540368 69018 540424
rect 69074 540368 71514 540424
rect 69013 540366 71514 540368
rect 69013 540363 69079 540366
rect 71454 540364 71514 540366
rect 71454 540304 72036 540364
rect 519892 538114 520474 538168
rect 522481 538114 522547 538117
rect 519892 538112 522547 538114
rect 519892 538108 522486 538112
rect 520414 538056 522486 538108
rect 522542 538056 522547 538112
rect 520414 538054 522547 538056
rect 522481 538051 522547 538054
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 69013 529274 69079 529277
rect 69013 529272 71514 529274
rect 69013 529216 69018 529272
rect 69074 529262 71514 529272
rect 69074 529216 72036 529262
rect 69013 529214 72036 529216
rect 69013 529211 69079 529214
rect 71454 529202 72036 529214
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 522297 515402 522363 515405
rect 520414 515400 522363 515402
rect 520414 515354 522302 515400
rect 519892 515344 522302 515354
rect 522358 515344 522363 515400
rect 519892 515342 522363 515344
rect 519892 515294 520474 515342
rect 522297 515339 522363 515342
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 69013 506970 69079 506973
rect 69013 506968 71514 506970
rect 69013 506912 69018 506968
rect 69074 506936 71514 506968
rect 69074 506912 72036 506936
rect 69013 506910 72036 506912
rect 69013 506907 69079 506910
rect 71454 506876 72036 506910
rect 519892 503978 520474 504008
rect 522389 503978 522455 503981
rect 519892 503976 522455 503978
rect 519892 503948 522394 503976
rect 520414 503920 522394 503948
rect 522450 503920 522455 503976
rect 520414 503918 522455 503920
rect 522389 503915 522455 503918
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect 69013 495682 69079 495685
rect 71454 495682 72036 495712
rect 69013 495680 72036 495682
rect 69013 495624 69018 495680
rect 69074 495652 72036 495680
rect 69074 495624 71514 495652
rect 69013 495622 71514 495624
rect 69013 495619 69079 495622
rect 522297 492554 522363 492557
rect 520414 492552 522363 492554
rect 520414 492540 522302 492552
rect 519892 492496 522302 492540
rect 522358 492496 522363 492552
rect 519892 492494 522363 492496
rect 519892 492480 520474 492494
rect 522297 492491 522363 492494
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 69013 484530 69079 484533
rect 69013 484528 71514 484530
rect 69013 484472 69018 484528
rect 69074 484488 71514 484528
rect 583520 484516 584960 484606
rect 69074 484472 72036 484488
rect 69013 484470 72036 484472
rect 69013 484467 69079 484470
rect 71454 484428 72036 484470
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 519892 469842 520474 469848
rect 522297 469842 522363 469845
rect 519892 469840 522363 469842
rect 519892 469788 522302 469840
rect 520414 469784 522302 469788
rect 522358 469784 522363 469840
rect 520414 469782 522363 469784
rect 522297 469779 522363 469782
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 69013 462226 69079 462229
rect 69013 462224 71514 462226
rect 69013 462168 69018 462224
rect 69074 462168 71514 462224
rect 69013 462166 71514 462168
rect 69013 462163 69079 462166
rect 71454 462162 71514 462166
rect 71454 462102 72036 462162
rect 522389 458418 522455 458421
rect 520414 458416 522455 458418
rect 520414 458380 522394 458416
rect 519892 458360 522394 458380
rect 522450 458360 522455 458416
rect 519892 458358 522455 458360
rect 519892 458320 520474 458358
rect 522389 458355 522455 458358
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 69013 451074 69079 451077
rect 69013 451072 71514 451074
rect 69013 451016 69018 451072
rect 69074 451060 71514 451072
rect 69074 451016 72036 451060
rect 69013 451014 72036 451016
rect 69013 451011 69079 451014
rect 71454 451000 72036 451014
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 519892 446994 520474 447034
rect 522297 446994 522363 446997
rect 519892 446992 522363 446994
rect 519892 446974 522302 446992
rect 520414 446936 522302 446974
rect 522358 446936 522363 446992
rect 520414 446934 522363 446936
rect 522297 446931 522363 446934
rect 583520 444668 584960 444908
rect 69013 439922 69079 439925
rect 69013 439920 71514 439922
rect 69013 439864 69018 439920
rect 69074 439864 71514 439920
rect 69013 439862 71514 439864
rect 69013 439859 69079 439862
rect 71454 439836 71514 439862
rect 71454 439776 72036 439836
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 522941 424282 523007 424285
rect 520414 424280 523007 424282
rect 520414 424224 522946 424280
rect 523002 424224 523007 424280
rect 520414 424222 523007 424224
rect 520414 424220 520474 424222
rect 519892 424160 520474 424220
rect 522941 424219 523007 424222
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 69013 417482 69079 417485
rect 71454 417482 72036 417510
rect 69013 417480 72036 417482
rect 69013 417424 69018 417480
rect 69074 417450 72036 417480
rect 69074 417424 71514 417450
rect 69013 417422 71514 417424
rect 69013 417419 69079 417422
rect 519892 412858 520474 412874
rect 522941 412858 523007 412861
rect 519892 412856 523007 412858
rect 519892 412814 522946 412856
rect 520414 412800 522946 412814
rect 523002 412800 523007 412856
rect 520414 412798 523007 412800
rect 522941 412795 523007 412798
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 69013 406466 69079 406469
rect 69013 406464 71514 406466
rect 69013 406408 69018 406464
rect 69074 406408 71514 406464
rect 69013 406406 72036 406408
rect 69013 406403 69079 406406
rect 71454 406348 72036 406406
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 522021 401570 522087 401573
rect 520414 401568 522087 401570
rect 520414 401528 522026 401568
rect 519892 401512 522026 401528
rect 522082 401512 522087 401568
rect 519892 401510 522087 401512
rect 519892 401468 520474 401510
rect 522021 401507 522087 401510
rect -960 397490 480 397580
rect 2865 397490 2931 397493
rect -960 397488 2931 397490
rect -960 397432 2870 397488
rect 2926 397432 2931 397488
rect -960 397430 2931 397432
rect -960 397340 480 397430
rect 2865 397427 2931 397430
rect 69013 395178 69079 395181
rect 71454 395178 72036 395184
rect 69013 395176 72036 395178
rect 69013 395120 69018 395176
rect 69074 395124 72036 395176
rect 69074 395120 71514 395124
rect 69013 395118 71514 395120
rect 69013 395115 69079 395118
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 522941 378722 523007 378725
rect 520414 378720 523007 378722
rect 520414 378714 522946 378720
rect 519892 378664 522946 378714
rect 523002 378664 523007 378720
rect 519892 378662 523007 378664
rect 519892 378654 520474 378662
rect 522941 378659 523007 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 69013 372874 69079 372877
rect 69013 372872 71514 372874
rect 69013 372816 69018 372872
rect 69074 372858 71514 372872
rect 69074 372816 72036 372858
rect 69013 372814 72036 372816
rect 69013 372811 69079 372814
rect 71454 372798 72036 372814
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 519892 367308 520474 367368
rect 520414 367298 520474 367308
rect 522941 367298 523007 367301
rect 520414 367296 523007 367298
rect 520414 367240 522946 367296
rect 523002 367240 523007 367296
rect 520414 367238 523007 367240
rect 522941 367235 523007 367238
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 69013 361722 69079 361725
rect 69013 361720 71514 361722
rect 69013 361664 69018 361720
rect 69074 361664 71514 361720
rect 69013 361662 71514 361664
rect 69013 361659 69079 361662
rect 71454 361634 71514 361662
rect 71454 361574 72036 361634
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 519892 356010 520474 356022
rect 522941 356010 523007 356013
rect 519892 356008 523007 356010
rect 519892 355962 522946 356008
rect 520414 355952 522946 355962
rect 523002 355952 523007 356008
rect 520414 355950 523007 355952
rect 522941 355947 523007 355950
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 71454 350472 72036 350532
rect 69013 350434 69079 350437
rect 71454 350434 71514 350472
rect 69013 350432 71514 350434
rect 69013 350376 69018 350432
rect 69074 350376 71514 350432
rect 69013 350374 71514 350376
rect 69013 350371 69079 350374
rect -960 345402 480 345492
rect 2865 345402 2931 345405
rect -960 345400 2931 345402
rect -960 345344 2870 345400
rect 2926 345344 2931 345400
rect -960 345342 2931 345344
rect -960 345252 480 345342
rect 2865 345339 2931 345342
rect 583520 338452 584960 338692
rect 519892 333162 520474 333208
rect 522297 333162 522363 333165
rect 519892 333160 522363 333162
rect 519892 333148 522302 333160
rect 520414 333104 522302 333148
rect 522358 333104 522363 333160
rect 520414 333102 522363 333104
rect 522297 333099 522363 333102
rect -960 332196 480 332436
rect 71454 328146 72036 328206
rect 69013 328130 69079 328133
rect 71454 328130 71514 328146
rect 69013 328128 71514 328130
rect 69013 328072 69018 328128
rect 69074 328072 71514 328128
rect 69013 328070 71514 328072
rect 69013 328067 69079 328070
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 522297 321874 522363 321877
rect 520414 321872 522363 321874
rect 520414 321862 522302 321872
rect 519892 321816 522302 321862
rect 522358 321816 522363 321872
rect 519892 321814 522363 321816
rect 519892 321802 520474 321814
rect 522297 321811 522363 321814
rect -960 319290 480 319380
rect 2865 319290 2931 319293
rect -960 319288 2931 319290
rect -960 319232 2870 319288
rect 2926 319232 2931 319288
rect -960 319230 2931 319232
rect -960 319140 480 319230
rect 2865 319227 2931 319230
rect 69013 316978 69079 316981
rect 71454 316978 72036 316982
rect 69013 316976 72036 316978
rect 69013 316920 69018 316976
rect 69074 316922 72036 316976
rect 69074 316920 71514 316922
rect 69013 316918 71514 316920
rect 69013 316915 69079 316918
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 519892 310334 520474 310394
rect 520414 310314 520474 310334
rect 522297 310314 522363 310317
rect 520414 310312 522363 310314
rect 520414 310256 522302 310312
rect 522358 310256 522363 310312
rect 520414 310254 522363 310256
rect 522297 310251 522363 310254
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 69013 305826 69079 305829
rect 71454 305826 72036 305880
rect 69013 305824 72036 305826
rect 69013 305768 69018 305824
rect 69074 305820 72036 305824
rect 69074 305768 71514 305820
rect 69013 305766 71514 305768
rect 69013 305763 69079 305766
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 522389 287738 522455 287741
rect 520414 287736 522455 287738
rect 520414 287702 522394 287736
rect 519892 287680 522394 287702
rect 522450 287680 522455 287736
rect 519892 287678 522455 287680
rect 519892 287642 520474 287678
rect 522389 287675 522455 287678
rect 583520 285276 584960 285516
rect 69013 283386 69079 283389
rect 71454 283386 72036 283432
rect 69013 283384 72036 283386
rect 69013 283328 69018 283384
rect 69074 283372 72036 283384
rect 69074 283328 71514 283372
rect 69013 283326 71514 283328
rect 69013 283323 69079 283326
rect -960 279972 480 280212
rect 519892 276178 520474 276234
rect 522297 276178 522363 276181
rect 519892 276176 522363 276178
rect 519892 276174 522302 276176
rect 520414 276120 522302 276174
rect 522358 276120 522363 276176
rect 520414 276118 522363 276120
rect 522297 276115 522363 276118
rect 69013 272370 69079 272373
rect 69013 272368 71514 272370
rect 69013 272312 69018 272368
rect 69074 272330 71514 272368
rect 69074 272312 72036 272330
rect 69013 272310 72036 272312
rect 69013 272307 69079 272310
rect 71454 272270 72036 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 522389 264890 522455 264893
rect 520414 264888 522455 264890
rect 519892 264832 522394 264888
rect 522450 264832 522455 264888
rect 519892 264830 522455 264832
rect 519892 264828 520474 264830
rect 522389 264827 522455 264830
rect 69013 261082 69079 261085
rect 71454 261082 72036 261106
rect 69013 261080 72036 261082
rect 69013 261024 69018 261080
rect 69074 261046 72036 261080
rect 69074 261024 71514 261046
rect 69013 261022 71514 261024
rect 69013 261019 69079 261022
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 519892 253482 520474 253542
rect 520414 253466 520474 253482
rect 522297 253466 522363 253469
rect 520414 253464 522363 253466
rect 520414 253408 522302 253464
rect 522358 253408 522363 253464
rect 520414 253406 522363 253408
rect 522297 253403 522363 253406
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 519892 242042 520474 242074
rect 522389 242042 522455 242045
rect 519892 242040 522455 242042
rect 519892 242014 522394 242040
rect 520414 241984 522394 242014
rect 522450 241984 522455 242040
rect 520414 241982 522455 241984
rect 522389 241979 522455 241982
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 69013 238778 69079 238781
rect 71454 238778 72036 238780
rect 69013 238776 72036 238778
rect 69013 238720 69018 238776
rect 69074 238720 72036 238776
rect 69013 238718 71514 238720
rect 69013 238715 69079 238718
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 522297 230754 522363 230757
rect 520414 230752 522363 230754
rect 520414 230728 522302 230752
rect 519892 230696 522302 230728
rect 522358 230696 522363 230752
rect 519892 230694 522363 230696
rect 519892 230668 520474 230694
rect 522297 230691 522363 230694
rect -960 227884 480 228124
rect 69013 227626 69079 227629
rect 71454 227626 72036 227678
rect 69013 227624 72036 227626
rect 69013 227568 69018 227624
rect 69074 227618 72036 227624
rect 69074 227568 71514 227618
rect 69013 227566 71514 227568
rect 69013 227563 69079 227566
rect 519892 219330 520474 219382
rect 522481 219330 522547 219333
rect 519892 219328 522547 219330
rect 519892 219322 522486 219328
rect 520414 219272 522486 219322
rect 522542 219272 522547 219328
rect 520414 219270 522547 219272
rect 522481 219267 522547 219270
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 69013 216474 69079 216477
rect 69013 216472 71514 216474
rect 69013 216416 69018 216472
rect 69074 216454 71514 216472
rect 69074 216416 72036 216454
rect 69013 216414 72036 216416
rect 69013 216411 69079 216414
rect 71454 216394 72036 216414
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 519892 207906 520474 207914
rect 522389 207906 522455 207909
rect 519892 207904 522455 207906
rect 519892 207854 522394 207904
rect 520414 207848 522394 207854
rect 522450 207848 522455 207904
rect 520414 207846 522455 207848
rect 522389 207843 522455 207846
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 519892 196508 520474 196568
rect 520414 196482 520474 196508
rect 522297 196482 522363 196485
rect 520414 196480 522363 196482
rect 520414 196424 522302 196480
rect 522358 196424 522363 196480
rect 520414 196422 522363 196424
rect 522297 196419 522363 196422
rect 69013 194170 69079 194173
rect 69013 194168 71514 194170
rect 69013 194112 69018 194168
rect 69074 194128 71514 194168
rect 69074 194112 72036 194128
rect 69013 194110 72036 194112
rect 69013 194107 69079 194110
rect 71454 194068 72036 194110
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 519892 185194 520474 185222
rect 522481 185194 522547 185197
rect 519892 185192 522547 185194
rect 519892 185162 522486 185192
rect 520414 185136 522486 185162
rect 522542 185136 522547 185192
rect 520414 185134 522547 185136
rect 522481 185131 522547 185134
rect 69013 182882 69079 182885
rect 71454 182882 72036 182904
rect 69013 182880 72036 182882
rect 69013 182824 69018 182880
rect 69074 182844 72036 182880
rect 69074 182824 71514 182844
rect 69013 182822 71514 182824
rect 69013 182819 69079 182822
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 522389 173906 522455 173909
rect 520414 173904 522455 173906
rect 520414 173876 522394 173904
rect 519892 173848 522394 173876
rect 522450 173848 522455 173904
rect 519892 173846 522455 173848
rect 519892 173816 520474 173846
rect 522389 173843 522455 173846
rect 71454 171742 72036 171802
rect 69013 171730 69079 171733
rect 71454 171730 71514 171742
rect 69013 171728 71514 171730
rect 69013 171672 69018 171728
rect 69074 171672 71514 171728
rect 69013 171670 71514 171672
rect 69013 171667 69079 171670
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3601 162890 3667 162893
rect -960 162888 3667 162890
rect -960 162832 3606 162888
rect 3662 162832 3667 162888
rect -960 162830 3667 162832
rect -960 162740 480 162830
rect 3601 162827 3667 162830
rect 519892 162348 520474 162408
rect 520414 162346 520474 162348
rect 522297 162346 522363 162349
rect 520414 162344 522363 162346
rect 520414 162288 522302 162344
rect 522358 162288 522363 162344
rect 520414 162286 522363 162288
rect 522297 162283 522363 162286
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 519892 151058 520474 151062
rect 522573 151058 522639 151061
rect 519892 151056 522639 151058
rect 519892 151002 522578 151056
rect 520414 151000 522578 151002
rect 522634 151000 522639 151056
rect 520414 150998 522639 151000
rect 522573 150995 522639 150998
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 69013 149426 69079 149429
rect 71454 149426 72036 149476
rect 69013 149424 72036 149426
rect 69013 149368 69018 149424
rect 69074 149416 72036 149424
rect 69074 149368 71514 149416
rect 69013 149366 71514 149368
rect 69013 149363 69079 149366
rect 519892 139656 520474 139716
rect 520414 139634 520474 139656
rect 522481 139634 522547 139637
rect 520414 139632 522547 139634
rect 520414 139576 522486 139632
rect 522542 139576 522547 139632
rect 520414 139574 522547 139576
rect 522481 139571 522547 139574
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 69013 138274 69079 138277
rect 69013 138272 71514 138274
rect 69013 138216 69018 138272
rect 69074 138252 71514 138272
rect 69074 138216 72036 138252
rect 69013 138214 72036 138216
rect 69013 138211 69079 138214
rect 71454 138192 72036 138214
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 519892 128210 520474 128248
rect 522389 128210 522455 128213
rect 519892 128208 522455 128210
rect 519892 128188 522394 128208
rect 520414 128152 522394 128188
rect 522450 128152 522455 128208
rect 520414 128150 522455 128152
rect 522389 128147 522455 128150
rect 69013 127122 69079 127125
rect 71454 127122 72036 127150
rect 69013 127120 72036 127122
rect 69013 127064 69018 127120
rect 69074 127090 72036 127120
rect 69074 127064 71514 127090
rect 69013 127062 71514 127064
rect 69013 127059 69079 127062
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 522297 116922 522363 116925
rect 520414 116920 522363 116922
rect 520414 116902 522302 116920
rect 519892 116864 522302 116902
rect 522358 116864 522363 116920
rect 519892 116862 522363 116864
rect 519892 116842 520474 116862
rect 522297 116859 522363 116862
rect 71454 115866 72036 115926
rect 69013 115834 69079 115837
rect 71454 115834 71514 115866
rect 69013 115832 71514 115834
rect 69013 115776 69018 115832
rect 69074 115776 71514 115832
rect 69013 115774 71514 115776
rect 69013 115771 69079 115774
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3693 110666 3759 110669
rect -960 110664 3759 110666
rect -960 110608 3698 110664
rect 3754 110608 3759 110664
rect -960 110606 3759 110608
rect -960 110516 480 110606
rect 3693 110603 3759 110606
rect 519892 105498 520474 105556
rect 522665 105498 522731 105501
rect 519892 105496 522731 105498
rect 520414 105440 522670 105496
rect 522726 105440 522731 105496
rect 520414 105438 522731 105440
rect 522665 105435 522731 105438
rect 69013 104818 69079 104821
rect 71454 104818 72036 104824
rect 69013 104816 72036 104818
rect 69013 104760 69018 104816
rect 69074 104764 72036 104816
rect 69074 104760 71514 104764
rect 69013 104758 71514 104760
rect 69013 104755 69079 104758
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 519892 94074 520474 94088
rect 522573 94074 522639 94077
rect 519892 94072 522639 94074
rect 519892 94028 522578 94072
rect 520414 94016 522578 94028
rect 522634 94016 522639 94072
rect 520414 94014 522639 94016
rect 522573 94011 522639 94014
rect 71454 93540 72036 93600
rect 69013 93530 69079 93533
rect 71454 93530 71514 93540
rect 69013 93528 71514 93530
rect 69013 93472 69018 93528
rect 69074 93472 71514 93528
rect 69013 93470 71514 93472
rect 69013 93467 69079 93470
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 522481 82786 522547 82789
rect 520414 82784 522547 82786
rect 520414 82742 522486 82784
rect 519892 82728 522486 82742
rect 522542 82728 522547 82784
rect 519892 82726 522547 82728
rect 519892 82682 520474 82726
rect 522481 82723 522547 82726
rect 69013 82378 69079 82381
rect 69013 82376 71514 82378
rect 69013 82320 69018 82376
rect 69074 82320 72036 82376
rect 69013 82318 72036 82320
rect 69013 82315 69079 82318
rect 71454 82316 72036 82318
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 519892 71362 520474 71396
rect 522389 71362 522455 71365
rect 519892 71360 522455 71362
rect 519892 71336 522394 71360
rect 520414 71304 522394 71336
rect 522450 71304 522455 71360
rect 520414 71302 522455 71304
rect 522389 71299 522455 71302
rect 69013 71226 69079 71229
rect 71454 71226 72036 71274
rect 69013 71224 72036 71226
rect 69013 71168 69018 71224
rect 69074 71214 72036 71224
rect 69074 71168 71514 71214
rect 69013 71166 71514 71168
rect 69013 71163 69079 71166
rect 69013 61162 69079 61165
rect 69013 61160 71514 61162
rect 69013 61104 69018 61160
rect 69074 61148 71514 61160
rect 69074 61104 72036 61148
rect 69013 61102 72036 61104
rect 69013 61099 69079 61102
rect 71454 61088 72036 61102
rect 519892 60890 520474 60904
rect 522297 60890 522363 60893
rect 519892 60888 522363 60890
rect 519892 60844 522302 60888
rect 520414 60832 522302 60844
rect 522358 60832 522363 60888
rect 520414 60830 522363 60832
rect 522297 60827 522363 60830
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3785 58578 3851 58581
rect -960 58576 3851 58578
rect -960 58520 3790 58576
rect 3846 58520 3851 58576
rect -960 58518 3851 58520
rect -960 58428 480 58518
rect 3785 58515 3851 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 365805 3770 365871 3773
rect 460933 3770 460999 3773
rect 365805 3768 460999 3770
rect 365805 3712 365810 3768
rect 365866 3712 460938 3768
rect 460994 3712 460999 3768
rect 365805 3710 460999 3712
rect 365805 3707 365871 3710
rect 460933 3707 460999 3710
rect 362309 3634 362375 3637
rect 459737 3634 459803 3637
rect 362309 3632 459803 3634
rect 362309 3576 362314 3632
rect 362370 3576 459742 3632
rect 459798 3576 459803 3632
rect 362309 3574 459803 3576
rect 362309 3571 362375 3574
rect 459737 3571 459803 3574
rect 358721 3498 358787 3501
rect 459645 3498 459711 3501
rect 358721 3496 459711 3498
rect 358721 3440 358726 3496
rect 358782 3440 459650 3496
rect 459706 3440 459711 3496
rect 358721 3438 459711 3440
rect 358721 3435 358787 3438
rect 459645 3435 459711 3438
rect 460933 3498 460999 3501
rect 462589 3498 462655 3501
rect 460933 3496 462655 3498
rect 460933 3440 460938 3496
rect 460994 3440 462594 3496
rect 462650 3440 462655 3496
rect 460933 3438 462655 3440
rect 460933 3435 460999 3438
rect 462589 3435 462655 3438
rect 355225 3362 355291 3365
rect 458173 3362 458239 3365
rect 355225 3360 458239 3362
rect 355225 3304 355230 3360
rect 355286 3304 458178 3360
rect 458234 3304 458239 3360
rect 355225 3302 458239 3304
rect 355225 3299 355291 3302
rect 458173 3299 458239 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 654008 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 654008 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 654008 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 654008 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 654008 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 654008 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 654008 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 654008 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 654008 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 654008 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 654008 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 654008 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 654008 128414 668898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 654008 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 654008 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 654008 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 654008 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 654008 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 654008 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 654008 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 654008 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 654008 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 654008 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 654008 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 654008 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 654008 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 654008 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 654008 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 654008 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 654008 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 654008 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 654008 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 654008 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 654008 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 654008 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 654008 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 654008 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 654008 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 654008 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 654008 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 654008 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 654008 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 654008 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 654008 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 654008 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 654008 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 654008 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 654008 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 654008 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 654008 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 654008 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 654008 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 654008 308414 668898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 654008 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 654008 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 654008 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 654008 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 654008 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 654008 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 654008 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 654008 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 654008 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 654008 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 654008 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 654008 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 654008 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 654008 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 654008 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 654008 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 654008 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 654008 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 654008 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 654008 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 654008 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 654008 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 654008 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 654008 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 654008 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 654008 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 654008 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 654008 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 654008 438134 654618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 654008 441854 658338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 654008 445574 662058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 654008 452414 668898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 654008 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 654008 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 654008 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 654008 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 654008 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 654008 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 654008 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 654008 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 654008 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 654008 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 654008 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 654008 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 654008 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 654008 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 654008 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 72798 633454 73798 633486
rect 72798 633218 72860 633454
rect 73096 633218 73180 633454
rect 73416 633218 73500 633454
rect 73736 633218 73798 633454
rect 72798 633134 73798 633218
rect 72798 632898 72860 633134
rect 73096 632898 73180 633134
rect 73416 632898 73500 633134
rect 73736 632898 73798 633134
rect 72798 632866 73798 632898
rect 518150 633454 519150 633486
rect 518150 633218 518212 633454
rect 518448 633218 518532 633454
rect 518768 633218 518852 633454
rect 519088 633218 519150 633454
rect 518150 633134 519150 633218
rect 518150 632898 518212 633134
rect 518448 632898 518532 633134
rect 518768 632898 518852 633134
rect 519088 632898 519150 633134
rect 518150 632866 519150 632898
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 74158 615454 75158 615486
rect 74158 615218 74220 615454
rect 74456 615218 74540 615454
rect 74776 615218 74860 615454
rect 75096 615218 75158 615454
rect 74158 615134 75158 615218
rect 74158 614898 74220 615134
rect 74456 614898 74540 615134
rect 74776 614898 74860 615134
rect 75096 614898 75158 615134
rect 74158 614866 75158 614898
rect 516790 615454 517790 615486
rect 516790 615218 516852 615454
rect 517088 615218 517172 615454
rect 517408 615218 517492 615454
rect 517728 615218 517790 615454
rect 516790 615134 517790 615218
rect 516790 614898 516852 615134
rect 517088 614898 517172 615134
rect 517408 614898 517492 615134
rect 517728 614898 517790 615134
rect 516790 614866 517790 614898
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 72798 597454 73798 597486
rect 72798 597218 72860 597454
rect 73096 597218 73180 597454
rect 73416 597218 73500 597454
rect 73736 597218 73798 597454
rect 72798 597134 73798 597218
rect 72798 596898 72860 597134
rect 73096 596898 73180 597134
rect 73416 596898 73500 597134
rect 73736 596898 73798 597134
rect 72798 596866 73798 596898
rect 518150 597454 519150 597486
rect 518150 597218 518212 597454
rect 518448 597218 518532 597454
rect 518768 597218 518852 597454
rect 519088 597218 519150 597454
rect 518150 597134 519150 597218
rect 518150 596898 518212 597134
rect 518448 596898 518532 597134
rect 518768 596898 518852 597134
rect 519088 596898 519150 597134
rect 518150 596866 519150 596898
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 74158 579454 75158 579486
rect 74158 579218 74220 579454
rect 74456 579218 74540 579454
rect 74776 579218 74860 579454
rect 75096 579218 75158 579454
rect 74158 579134 75158 579218
rect 74158 578898 74220 579134
rect 74456 578898 74540 579134
rect 74776 578898 74860 579134
rect 75096 578898 75158 579134
rect 74158 578866 75158 578898
rect 516790 579454 517790 579486
rect 516790 579218 516852 579454
rect 517088 579218 517172 579454
rect 517408 579218 517492 579454
rect 517728 579218 517790 579454
rect 516790 579134 517790 579218
rect 516790 578898 516852 579134
rect 517088 578898 517172 579134
rect 517408 578898 517492 579134
rect 517728 578898 517790 579134
rect 516790 578866 517790 578898
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 72798 561454 73798 561486
rect 72798 561218 72860 561454
rect 73096 561218 73180 561454
rect 73416 561218 73500 561454
rect 73736 561218 73798 561454
rect 72798 561134 73798 561218
rect 72798 560898 72860 561134
rect 73096 560898 73180 561134
rect 73416 560898 73500 561134
rect 73736 560898 73798 561134
rect 72798 560866 73798 560898
rect 518150 561454 519150 561486
rect 518150 561218 518212 561454
rect 518448 561218 518532 561454
rect 518768 561218 518852 561454
rect 519088 561218 519150 561454
rect 518150 561134 519150 561218
rect 518150 560898 518212 561134
rect 518448 560898 518532 561134
rect 518768 560898 518852 561134
rect 519088 560898 519150 561134
rect 518150 560866 519150 560898
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 74158 543454 75158 543486
rect 74158 543218 74220 543454
rect 74456 543218 74540 543454
rect 74776 543218 74860 543454
rect 75096 543218 75158 543454
rect 74158 543134 75158 543218
rect 74158 542898 74220 543134
rect 74456 542898 74540 543134
rect 74776 542898 74860 543134
rect 75096 542898 75158 543134
rect 74158 542866 75158 542898
rect 516790 543454 517790 543486
rect 516790 543218 516852 543454
rect 517088 543218 517172 543454
rect 517408 543218 517492 543454
rect 517728 543218 517790 543454
rect 516790 543134 517790 543218
rect 516790 542898 516852 543134
rect 517088 542898 517172 543134
rect 517408 542898 517492 543134
rect 517728 542898 517790 543134
rect 516790 542866 517790 542898
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 72798 525454 73798 525486
rect 72798 525218 72860 525454
rect 73096 525218 73180 525454
rect 73416 525218 73500 525454
rect 73736 525218 73798 525454
rect 72798 525134 73798 525218
rect 72798 524898 72860 525134
rect 73096 524898 73180 525134
rect 73416 524898 73500 525134
rect 73736 524898 73798 525134
rect 72798 524866 73798 524898
rect 518150 525454 519150 525486
rect 518150 525218 518212 525454
rect 518448 525218 518532 525454
rect 518768 525218 518852 525454
rect 519088 525218 519150 525454
rect 518150 525134 519150 525218
rect 518150 524898 518212 525134
rect 518448 524898 518532 525134
rect 518768 524898 518852 525134
rect 519088 524898 519150 525134
rect 518150 524866 519150 524898
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 74158 507454 75158 507486
rect 74158 507218 74220 507454
rect 74456 507218 74540 507454
rect 74776 507218 74860 507454
rect 75096 507218 75158 507454
rect 74158 507134 75158 507218
rect 74158 506898 74220 507134
rect 74456 506898 74540 507134
rect 74776 506898 74860 507134
rect 75096 506898 75158 507134
rect 74158 506866 75158 506898
rect 516790 507454 517790 507486
rect 516790 507218 516852 507454
rect 517088 507218 517172 507454
rect 517408 507218 517492 507454
rect 517728 507218 517790 507454
rect 516790 507134 517790 507218
rect 516790 506898 516852 507134
rect 517088 506898 517172 507134
rect 517408 506898 517492 507134
rect 517728 506898 517790 507134
rect 516790 506866 517790 506898
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 72798 489454 73798 489486
rect 72798 489218 72860 489454
rect 73096 489218 73180 489454
rect 73416 489218 73500 489454
rect 73736 489218 73798 489454
rect 72798 489134 73798 489218
rect 72798 488898 72860 489134
rect 73096 488898 73180 489134
rect 73416 488898 73500 489134
rect 73736 488898 73798 489134
rect 72798 488866 73798 488898
rect 518150 489454 519150 489486
rect 518150 489218 518212 489454
rect 518448 489218 518532 489454
rect 518768 489218 518852 489454
rect 519088 489218 519150 489454
rect 518150 489134 519150 489218
rect 518150 488898 518212 489134
rect 518448 488898 518532 489134
rect 518768 488898 518852 489134
rect 519088 488898 519150 489134
rect 518150 488866 519150 488898
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 74158 471454 75158 471486
rect 74158 471218 74220 471454
rect 74456 471218 74540 471454
rect 74776 471218 74860 471454
rect 75096 471218 75158 471454
rect 74158 471134 75158 471218
rect 74158 470898 74220 471134
rect 74456 470898 74540 471134
rect 74776 470898 74860 471134
rect 75096 470898 75158 471134
rect 74158 470866 75158 470898
rect 516790 471454 517790 471486
rect 516790 471218 516852 471454
rect 517088 471218 517172 471454
rect 517408 471218 517492 471454
rect 517728 471218 517790 471454
rect 516790 471134 517790 471218
rect 516790 470898 516852 471134
rect 517088 470898 517172 471134
rect 517408 470898 517492 471134
rect 517728 470898 517790 471134
rect 516790 470866 517790 470898
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 72798 453454 73798 453486
rect 72798 453218 72860 453454
rect 73096 453218 73180 453454
rect 73416 453218 73500 453454
rect 73736 453218 73798 453454
rect 72798 453134 73798 453218
rect 72798 452898 72860 453134
rect 73096 452898 73180 453134
rect 73416 452898 73500 453134
rect 73736 452898 73798 453134
rect 72798 452866 73798 452898
rect 518150 453454 519150 453486
rect 518150 453218 518212 453454
rect 518448 453218 518532 453454
rect 518768 453218 518852 453454
rect 519088 453218 519150 453454
rect 518150 453134 519150 453218
rect 518150 452898 518212 453134
rect 518448 452898 518532 453134
rect 518768 452898 518852 453134
rect 519088 452898 519150 453134
rect 518150 452866 519150 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 74158 435454 75158 435486
rect 74158 435218 74220 435454
rect 74456 435218 74540 435454
rect 74776 435218 74860 435454
rect 75096 435218 75158 435454
rect 74158 435134 75158 435218
rect 74158 434898 74220 435134
rect 74456 434898 74540 435134
rect 74776 434898 74860 435134
rect 75096 434898 75158 435134
rect 74158 434866 75158 434898
rect 516790 435454 517790 435486
rect 516790 435218 516852 435454
rect 517088 435218 517172 435454
rect 517408 435218 517492 435454
rect 517728 435218 517790 435454
rect 516790 435134 517790 435218
rect 516790 434898 516852 435134
rect 517088 434898 517172 435134
rect 517408 434898 517492 435134
rect 517728 434898 517790 435134
rect 516790 434866 517790 434898
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 72798 417454 73798 417486
rect 72798 417218 72860 417454
rect 73096 417218 73180 417454
rect 73416 417218 73500 417454
rect 73736 417218 73798 417454
rect 72798 417134 73798 417218
rect 72798 416898 72860 417134
rect 73096 416898 73180 417134
rect 73416 416898 73500 417134
rect 73736 416898 73798 417134
rect 72798 416866 73798 416898
rect 518150 417454 519150 417486
rect 518150 417218 518212 417454
rect 518448 417218 518532 417454
rect 518768 417218 518852 417454
rect 519088 417218 519150 417454
rect 518150 417134 519150 417218
rect 518150 416898 518212 417134
rect 518448 416898 518532 417134
rect 518768 416898 518852 417134
rect 519088 416898 519150 417134
rect 518150 416866 519150 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 74158 399454 75158 399486
rect 74158 399218 74220 399454
rect 74456 399218 74540 399454
rect 74776 399218 74860 399454
rect 75096 399218 75158 399454
rect 74158 399134 75158 399218
rect 74158 398898 74220 399134
rect 74456 398898 74540 399134
rect 74776 398898 74860 399134
rect 75096 398898 75158 399134
rect 74158 398866 75158 398898
rect 516790 399454 517790 399486
rect 516790 399218 516852 399454
rect 517088 399218 517172 399454
rect 517408 399218 517492 399454
rect 517728 399218 517790 399454
rect 516790 399134 517790 399218
rect 516790 398898 516852 399134
rect 517088 398898 517172 399134
rect 517408 398898 517492 399134
rect 517728 398898 517790 399134
rect 516790 398866 517790 398898
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 72798 381454 73798 381486
rect 72798 381218 72860 381454
rect 73096 381218 73180 381454
rect 73416 381218 73500 381454
rect 73736 381218 73798 381454
rect 72798 381134 73798 381218
rect 72798 380898 72860 381134
rect 73096 380898 73180 381134
rect 73416 380898 73500 381134
rect 73736 380898 73798 381134
rect 72798 380866 73798 380898
rect 518150 381454 519150 381486
rect 518150 381218 518212 381454
rect 518448 381218 518532 381454
rect 518768 381218 518852 381454
rect 519088 381218 519150 381454
rect 518150 381134 519150 381218
rect 518150 380898 518212 381134
rect 518448 380898 518532 381134
rect 518768 380898 518852 381134
rect 519088 380898 519150 381134
rect 518150 380866 519150 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 74158 363454 75158 363486
rect 74158 363218 74220 363454
rect 74456 363218 74540 363454
rect 74776 363218 74860 363454
rect 75096 363218 75158 363454
rect 74158 363134 75158 363218
rect 74158 362898 74220 363134
rect 74456 362898 74540 363134
rect 74776 362898 74860 363134
rect 75096 362898 75158 363134
rect 74158 362866 75158 362898
rect 516790 363454 517790 363486
rect 516790 363218 516852 363454
rect 517088 363218 517172 363454
rect 517408 363218 517492 363454
rect 517728 363218 517790 363454
rect 516790 363134 517790 363218
rect 516790 362898 516852 363134
rect 517088 362898 517172 363134
rect 517408 362898 517492 363134
rect 517728 362898 517790 363134
rect 516790 362866 517790 362898
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 72798 345454 73798 345486
rect 72798 345218 72860 345454
rect 73096 345218 73180 345454
rect 73416 345218 73500 345454
rect 73736 345218 73798 345454
rect 72798 345134 73798 345218
rect 72798 344898 72860 345134
rect 73096 344898 73180 345134
rect 73416 344898 73500 345134
rect 73736 344898 73798 345134
rect 72798 344866 73798 344898
rect 518150 345454 519150 345486
rect 518150 345218 518212 345454
rect 518448 345218 518532 345454
rect 518768 345218 518852 345454
rect 519088 345218 519150 345454
rect 518150 345134 519150 345218
rect 518150 344898 518212 345134
rect 518448 344898 518532 345134
rect 518768 344898 518852 345134
rect 519088 344898 519150 345134
rect 518150 344866 519150 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 74158 327454 75158 327486
rect 74158 327218 74220 327454
rect 74456 327218 74540 327454
rect 74776 327218 74860 327454
rect 75096 327218 75158 327454
rect 74158 327134 75158 327218
rect 74158 326898 74220 327134
rect 74456 326898 74540 327134
rect 74776 326898 74860 327134
rect 75096 326898 75158 327134
rect 74158 326866 75158 326898
rect 516790 327454 517790 327486
rect 516790 327218 516852 327454
rect 517088 327218 517172 327454
rect 517408 327218 517492 327454
rect 517728 327218 517790 327454
rect 516790 327134 517790 327218
rect 516790 326898 516852 327134
rect 517088 326898 517172 327134
rect 517408 326898 517492 327134
rect 517728 326898 517790 327134
rect 516790 326866 517790 326898
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 72798 309454 73798 309486
rect 72798 309218 72860 309454
rect 73096 309218 73180 309454
rect 73416 309218 73500 309454
rect 73736 309218 73798 309454
rect 72798 309134 73798 309218
rect 72798 308898 72860 309134
rect 73096 308898 73180 309134
rect 73416 308898 73500 309134
rect 73736 308898 73798 309134
rect 72798 308866 73798 308898
rect 518150 309454 519150 309486
rect 518150 309218 518212 309454
rect 518448 309218 518532 309454
rect 518768 309218 518852 309454
rect 519088 309218 519150 309454
rect 518150 309134 519150 309218
rect 518150 308898 518212 309134
rect 518448 308898 518532 309134
rect 518768 308898 518852 309134
rect 519088 308898 519150 309134
rect 518150 308866 519150 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 74158 291454 75158 291486
rect 74158 291218 74220 291454
rect 74456 291218 74540 291454
rect 74776 291218 74860 291454
rect 75096 291218 75158 291454
rect 74158 291134 75158 291218
rect 74158 290898 74220 291134
rect 74456 290898 74540 291134
rect 74776 290898 74860 291134
rect 75096 290898 75158 291134
rect 74158 290866 75158 290898
rect 516790 291454 517790 291486
rect 516790 291218 516852 291454
rect 517088 291218 517172 291454
rect 517408 291218 517492 291454
rect 517728 291218 517790 291454
rect 516790 291134 517790 291218
rect 516790 290898 516852 291134
rect 517088 290898 517172 291134
rect 517408 290898 517492 291134
rect 517728 290898 517790 291134
rect 516790 290866 517790 290898
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 72798 273454 73798 273486
rect 72798 273218 72860 273454
rect 73096 273218 73180 273454
rect 73416 273218 73500 273454
rect 73736 273218 73798 273454
rect 72798 273134 73798 273218
rect 72798 272898 72860 273134
rect 73096 272898 73180 273134
rect 73416 272898 73500 273134
rect 73736 272898 73798 273134
rect 72798 272866 73798 272898
rect 518150 273454 519150 273486
rect 518150 273218 518212 273454
rect 518448 273218 518532 273454
rect 518768 273218 518852 273454
rect 519088 273218 519150 273454
rect 518150 273134 519150 273218
rect 518150 272898 518212 273134
rect 518448 272898 518532 273134
rect 518768 272898 518852 273134
rect 519088 272898 519150 273134
rect 518150 272866 519150 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 74158 255454 75158 255486
rect 74158 255218 74220 255454
rect 74456 255218 74540 255454
rect 74776 255218 74860 255454
rect 75096 255218 75158 255454
rect 74158 255134 75158 255218
rect 74158 254898 74220 255134
rect 74456 254898 74540 255134
rect 74776 254898 74860 255134
rect 75096 254898 75158 255134
rect 74158 254866 75158 254898
rect 516790 255454 517790 255486
rect 516790 255218 516852 255454
rect 517088 255218 517172 255454
rect 517408 255218 517492 255454
rect 517728 255218 517790 255454
rect 516790 255134 517790 255218
rect 516790 254898 516852 255134
rect 517088 254898 517172 255134
rect 517408 254898 517492 255134
rect 517728 254898 517790 255134
rect 516790 254866 517790 254898
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 72798 237454 73798 237486
rect 72798 237218 72860 237454
rect 73096 237218 73180 237454
rect 73416 237218 73500 237454
rect 73736 237218 73798 237454
rect 72798 237134 73798 237218
rect 72798 236898 72860 237134
rect 73096 236898 73180 237134
rect 73416 236898 73500 237134
rect 73736 236898 73798 237134
rect 72798 236866 73798 236898
rect 518150 237454 519150 237486
rect 518150 237218 518212 237454
rect 518448 237218 518532 237454
rect 518768 237218 518852 237454
rect 519088 237218 519150 237454
rect 518150 237134 519150 237218
rect 518150 236898 518212 237134
rect 518448 236898 518532 237134
rect 518768 236898 518852 237134
rect 519088 236898 519150 237134
rect 518150 236866 519150 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 74158 219454 75158 219486
rect 74158 219218 74220 219454
rect 74456 219218 74540 219454
rect 74776 219218 74860 219454
rect 75096 219218 75158 219454
rect 74158 219134 75158 219218
rect 74158 218898 74220 219134
rect 74456 218898 74540 219134
rect 74776 218898 74860 219134
rect 75096 218898 75158 219134
rect 74158 218866 75158 218898
rect 516790 219454 517790 219486
rect 516790 219218 516852 219454
rect 517088 219218 517172 219454
rect 517408 219218 517492 219454
rect 517728 219218 517790 219454
rect 516790 219134 517790 219218
rect 516790 218898 516852 219134
rect 517088 218898 517172 219134
rect 517408 218898 517492 219134
rect 517728 218898 517790 219134
rect 516790 218866 517790 218898
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 72798 201454 73798 201486
rect 72798 201218 72860 201454
rect 73096 201218 73180 201454
rect 73416 201218 73500 201454
rect 73736 201218 73798 201454
rect 72798 201134 73798 201218
rect 72798 200898 72860 201134
rect 73096 200898 73180 201134
rect 73416 200898 73500 201134
rect 73736 200898 73798 201134
rect 72798 200866 73798 200898
rect 518150 201454 519150 201486
rect 518150 201218 518212 201454
rect 518448 201218 518532 201454
rect 518768 201218 518852 201454
rect 519088 201218 519150 201454
rect 518150 201134 519150 201218
rect 518150 200898 518212 201134
rect 518448 200898 518532 201134
rect 518768 200898 518852 201134
rect 519088 200898 519150 201134
rect 518150 200866 519150 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 74158 183454 75158 183486
rect 74158 183218 74220 183454
rect 74456 183218 74540 183454
rect 74776 183218 74860 183454
rect 75096 183218 75158 183454
rect 74158 183134 75158 183218
rect 74158 182898 74220 183134
rect 74456 182898 74540 183134
rect 74776 182898 74860 183134
rect 75096 182898 75158 183134
rect 74158 182866 75158 182898
rect 516790 183454 517790 183486
rect 516790 183218 516852 183454
rect 517088 183218 517172 183454
rect 517408 183218 517492 183454
rect 517728 183218 517790 183454
rect 516790 183134 517790 183218
rect 516790 182898 516852 183134
rect 517088 182898 517172 183134
rect 517408 182898 517492 183134
rect 517728 182898 517790 183134
rect 516790 182866 517790 182898
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 72798 165454 73798 165486
rect 72798 165218 72860 165454
rect 73096 165218 73180 165454
rect 73416 165218 73500 165454
rect 73736 165218 73798 165454
rect 72798 165134 73798 165218
rect 72798 164898 72860 165134
rect 73096 164898 73180 165134
rect 73416 164898 73500 165134
rect 73736 164898 73798 165134
rect 72798 164866 73798 164898
rect 518150 165454 519150 165486
rect 518150 165218 518212 165454
rect 518448 165218 518532 165454
rect 518768 165218 518852 165454
rect 519088 165218 519150 165454
rect 518150 165134 519150 165218
rect 518150 164898 518212 165134
rect 518448 164898 518532 165134
rect 518768 164898 518852 165134
rect 519088 164898 519150 165134
rect 518150 164866 519150 164898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 74158 147454 75158 147486
rect 74158 147218 74220 147454
rect 74456 147218 74540 147454
rect 74776 147218 74860 147454
rect 75096 147218 75158 147454
rect 74158 147134 75158 147218
rect 74158 146898 74220 147134
rect 74456 146898 74540 147134
rect 74776 146898 74860 147134
rect 75096 146898 75158 147134
rect 74158 146866 75158 146898
rect 516790 147454 517790 147486
rect 516790 147218 516852 147454
rect 517088 147218 517172 147454
rect 517408 147218 517492 147454
rect 517728 147218 517790 147454
rect 516790 147134 517790 147218
rect 516790 146898 516852 147134
rect 517088 146898 517172 147134
rect 517408 146898 517492 147134
rect 517728 146898 517790 147134
rect 516790 146866 517790 146898
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 72798 129454 73798 129486
rect 72798 129218 72860 129454
rect 73096 129218 73180 129454
rect 73416 129218 73500 129454
rect 73736 129218 73798 129454
rect 72798 129134 73798 129218
rect 72798 128898 72860 129134
rect 73096 128898 73180 129134
rect 73416 128898 73500 129134
rect 73736 128898 73798 129134
rect 72798 128866 73798 128898
rect 518150 129454 519150 129486
rect 518150 129218 518212 129454
rect 518448 129218 518532 129454
rect 518768 129218 518852 129454
rect 519088 129218 519150 129454
rect 518150 129134 519150 129218
rect 518150 128898 518212 129134
rect 518448 128898 518532 129134
rect 518768 128898 518852 129134
rect 519088 128898 519150 129134
rect 518150 128866 519150 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 74158 111454 75158 111486
rect 74158 111218 74220 111454
rect 74456 111218 74540 111454
rect 74776 111218 74860 111454
rect 75096 111218 75158 111454
rect 74158 111134 75158 111218
rect 74158 110898 74220 111134
rect 74456 110898 74540 111134
rect 74776 110898 74860 111134
rect 75096 110898 75158 111134
rect 74158 110866 75158 110898
rect 516790 111454 517790 111486
rect 516790 111218 516852 111454
rect 517088 111218 517172 111454
rect 517408 111218 517492 111454
rect 517728 111218 517790 111454
rect 516790 111134 517790 111218
rect 516790 110898 516852 111134
rect 517088 110898 517172 111134
rect 517408 110898 517492 111134
rect 517728 110898 517790 111134
rect 516790 110866 517790 110898
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 72798 93454 73798 93486
rect 72798 93218 72860 93454
rect 73096 93218 73180 93454
rect 73416 93218 73500 93454
rect 73736 93218 73798 93454
rect 72798 93134 73798 93218
rect 72798 92898 72860 93134
rect 73096 92898 73180 93134
rect 73416 92898 73500 93134
rect 73736 92898 73798 93134
rect 72798 92866 73798 92898
rect 518150 93454 519150 93486
rect 518150 93218 518212 93454
rect 518448 93218 518532 93454
rect 518768 93218 518852 93454
rect 519088 93218 519150 93454
rect 518150 93134 519150 93218
rect 518150 92898 518212 93134
rect 518448 92898 518532 93134
rect 518768 92898 518852 93134
rect 519088 92898 519150 93134
rect 518150 92866 519150 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 74158 75454 75158 75486
rect 74158 75218 74220 75454
rect 74456 75218 74540 75454
rect 74776 75218 74860 75454
rect 75096 75218 75158 75454
rect 74158 75134 75158 75218
rect 74158 74898 74220 75134
rect 74456 74898 74540 75134
rect 74776 74898 74860 75134
rect 75096 74898 75158 75134
rect 74158 74866 75158 74898
rect 516790 75454 517790 75486
rect 516790 75218 516852 75454
rect 517088 75218 517172 75454
rect 517408 75218 517492 75454
rect 517728 75218 517790 75454
rect 516790 75134 517790 75218
rect 516790 74898 516852 75134
rect 517088 74898 517172 75134
rect 517408 74898 517492 75134
rect 517728 74898 517790 75134
rect 516790 74866 517790 74898
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 72860 633218 73096 633454
rect 73180 633218 73416 633454
rect 73500 633218 73736 633454
rect 72860 632898 73096 633134
rect 73180 632898 73416 633134
rect 73500 632898 73736 633134
rect 518212 633218 518448 633454
rect 518532 633218 518768 633454
rect 518852 633218 519088 633454
rect 518212 632898 518448 633134
rect 518532 632898 518768 633134
rect 518852 632898 519088 633134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 74220 615218 74456 615454
rect 74540 615218 74776 615454
rect 74860 615218 75096 615454
rect 74220 614898 74456 615134
rect 74540 614898 74776 615134
rect 74860 614898 75096 615134
rect 516852 615218 517088 615454
rect 517172 615218 517408 615454
rect 517492 615218 517728 615454
rect 516852 614898 517088 615134
rect 517172 614898 517408 615134
rect 517492 614898 517728 615134
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 72860 597218 73096 597454
rect 73180 597218 73416 597454
rect 73500 597218 73736 597454
rect 72860 596898 73096 597134
rect 73180 596898 73416 597134
rect 73500 596898 73736 597134
rect 518212 597218 518448 597454
rect 518532 597218 518768 597454
rect 518852 597218 519088 597454
rect 518212 596898 518448 597134
rect 518532 596898 518768 597134
rect 518852 596898 519088 597134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 74220 579218 74456 579454
rect 74540 579218 74776 579454
rect 74860 579218 75096 579454
rect 74220 578898 74456 579134
rect 74540 578898 74776 579134
rect 74860 578898 75096 579134
rect 516852 579218 517088 579454
rect 517172 579218 517408 579454
rect 517492 579218 517728 579454
rect 516852 578898 517088 579134
rect 517172 578898 517408 579134
rect 517492 578898 517728 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 72860 561218 73096 561454
rect 73180 561218 73416 561454
rect 73500 561218 73736 561454
rect 72860 560898 73096 561134
rect 73180 560898 73416 561134
rect 73500 560898 73736 561134
rect 518212 561218 518448 561454
rect 518532 561218 518768 561454
rect 518852 561218 519088 561454
rect 518212 560898 518448 561134
rect 518532 560898 518768 561134
rect 518852 560898 519088 561134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 74220 543218 74456 543454
rect 74540 543218 74776 543454
rect 74860 543218 75096 543454
rect 74220 542898 74456 543134
rect 74540 542898 74776 543134
rect 74860 542898 75096 543134
rect 516852 543218 517088 543454
rect 517172 543218 517408 543454
rect 517492 543218 517728 543454
rect 516852 542898 517088 543134
rect 517172 542898 517408 543134
rect 517492 542898 517728 543134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 72860 525218 73096 525454
rect 73180 525218 73416 525454
rect 73500 525218 73736 525454
rect 72860 524898 73096 525134
rect 73180 524898 73416 525134
rect 73500 524898 73736 525134
rect 518212 525218 518448 525454
rect 518532 525218 518768 525454
rect 518852 525218 519088 525454
rect 518212 524898 518448 525134
rect 518532 524898 518768 525134
rect 518852 524898 519088 525134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 74220 507218 74456 507454
rect 74540 507218 74776 507454
rect 74860 507218 75096 507454
rect 74220 506898 74456 507134
rect 74540 506898 74776 507134
rect 74860 506898 75096 507134
rect 516852 507218 517088 507454
rect 517172 507218 517408 507454
rect 517492 507218 517728 507454
rect 516852 506898 517088 507134
rect 517172 506898 517408 507134
rect 517492 506898 517728 507134
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 72860 489218 73096 489454
rect 73180 489218 73416 489454
rect 73500 489218 73736 489454
rect 72860 488898 73096 489134
rect 73180 488898 73416 489134
rect 73500 488898 73736 489134
rect 518212 489218 518448 489454
rect 518532 489218 518768 489454
rect 518852 489218 519088 489454
rect 518212 488898 518448 489134
rect 518532 488898 518768 489134
rect 518852 488898 519088 489134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 74220 471218 74456 471454
rect 74540 471218 74776 471454
rect 74860 471218 75096 471454
rect 74220 470898 74456 471134
rect 74540 470898 74776 471134
rect 74860 470898 75096 471134
rect 516852 471218 517088 471454
rect 517172 471218 517408 471454
rect 517492 471218 517728 471454
rect 516852 470898 517088 471134
rect 517172 470898 517408 471134
rect 517492 470898 517728 471134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 72860 453218 73096 453454
rect 73180 453218 73416 453454
rect 73500 453218 73736 453454
rect 72860 452898 73096 453134
rect 73180 452898 73416 453134
rect 73500 452898 73736 453134
rect 518212 453218 518448 453454
rect 518532 453218 518768 453454
rect 518852 453218 519088 453454
rect 518212 452898 518448 453134
rect 518532 452898 518768 453134
rect 518852 452898 519088 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 74220 435218 74456 435454
rect 74540 435218 74776 435454
rect 74860 435218 75096 435454
rect 74220 434898 74456 435134
rect 74540 434898 74776 435134
rect 74860 434898 75096 435134
rect 516852 435218 517088 435454
rect 517172 435218 517408 435454
rect 517492 435218 517728 435454
rect 516852 434898 517088 435134
rect 517172 434898 517408 435134
rect 517492 434898 517728 435134
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 72860 417218 73096 417454
rect 73180 417218 73416 417454
rect 73500 417218 73736 417454
rect 72860 416898 73096 417134
rect 73180 416898 73416 417134
rect 73500 416898 73736 417134
rect 518212 417218 518448 417454
rect 518532 417218 518768 417454
rect 518852 417218 519088 417454
rect 518212 416898 518448 417134
rect 518532 416898 518768 417134
rect 518852 416898 519088 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 74220 399218 74456 399454
rect 74540 399218 74776 399454
rect 74860 399218 75096 399454
rect 74220 398898 74456 399134
rect 74540 398898 74776 399134
rect 74860 398898 75096 399134
rect 516852 399218 517088 399454
rect 517172 399218 517408 399454
rect 517492 399218 517728 399454
rect 516852 398898 517088 399134
rect 517172 398898 517408 399134
rect 517492 398898 517728 399134
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 72860 381218 73096 381454
rect 73180 381218 73416 381454
rect 73500 381218 73736 381454
rect 72860 380898 73096 381134
rect 73180 380898 73416 381134
rect 73500 380898 73736 381134
rect 518212 381218 518448 381454
rect 518532 381218 518768 381454
rect 518852 381218 519088 381454
rect 518212 380898 518448 381134
rect 518532 380898 518768 381134
rect 518852 380898 519088 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 74220 363218 74456 363454
rect 74540 363218 74776 363454
rect 74860 363218 75096 363454
rect 74220 362898 74456 363134
rect 74540 362898 74776 363134
rect 74860 362898 75096 363134
rect 516852 363218 517088 363454
rect 517172 363218 517408 363454
rect 517492 363218 517728 363454
rect 516852 362898 517088 363134
rect 517172 362898 517408 363134
rect 517492 362898 517728 363134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 72860 345218 73096 345454
rect 73180 345218 73416 345454
rect 73500 345218 73736 345454
rect 72860 344898 73096 345134
rect 73180 344898 73416 345134
rect 73500 344898 73736 345134
rect 518212 345218 518448 345454
rect 518532 345218 518768 345454
rect 518852 345218 519088 345454
rect 518212 344898 518448 345134
rect 518532 344898 518768 345134
rect 518852 344898 519088 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 74220 327218 74456 327454
rect 74540 327218 74776 327454
rect 74860 327218 75096 327454
rect 74220 326898 74456 327134
rect 74540 326898 74776 327134
rect 74860 326898 75096 327134
rect 516852 327218 517088 327454
rect 517172 327218 517408 327454
rect 517492 327218 517728 327454
rect 516852 326898 517088 327134
rect 517172 326898 517408 327134
rect 517492 326898 517728 327134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 72860 309218 73096 309454
rect 73180 309218 73416 309454
rect 73500 309218 73736 309454
rect 72860 308898 73096 309134
rect 73180 308898 73416 309134
rect 73500 308898 73736 309134
rect 518212 309218 518448 309454
rect 518532 309218 518768 309454
rect 518852 309218 519088 309454
rect 518212 308898 518448 309134
rect 518532 308898 518768 309134
rect 518852 308898 519088 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 74220 291218 74456 291454
rect 74540 291218 74776 291454
rect 74860 291218 75096 291454
rect 74220 290898 74456 291134
rect 74540 290898 74776 291134
rect 74860 290898 75096 291134
rect 516852 291218 517088 291454
rect 517172 291218 517408 291454
rect 517492 291218 517728 291454
rect 516852 290898 517088 291134
rect 517172 290898 517408 291134
rect 517492 290898 517728 291134
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 72860 273218 73096 273454
rect 73180 273218 73416 273454
rect 73500 273218 73736 273454
rect 72860 272898 73096 273134
rect 73180 272898 73416 273134
rect 73500 272898 73736 273134
rect 518212 273218 518448 273454
rect 518532 273218 518768 273454
rect 518852 273218 519088 273454
rect 518212 272898 518448 273134
rect 518532 272898 518768 273134
rect 518852 272898 519088 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 74220 255218 74456 255454
rect 74540 255218 74776 255454
rect 74860 255218 75096 255454
rect 74220 254898 74456 255134
rect 74540 254898 74776 255134
rect 74860 254898 75096 255134
rect 516852 255218 517088 255454
rect 517172 255218 517408 255454
rect 517492 255218 517728 255454
rect 516852 254898 517088 255134
rect 517172 254898 517408 255134
rect 517492 254898 517728 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 72860 237218 73096 237454
rect 73180 237218 73416 237454
rect 73500 237218 73736 237454
rect 72860 236898 73096 237134
rect 73180 236898 73416 237134
rect 73500 236898 73736 237134
rect 518212 237218 518448 237454
rect 518532 237218 518768 237454
rect 518852 237218 519088 237454
rect 518212 236898 518448 237134
rect 518532 236898 518768 237134
rect 518852 236898 519088 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 74220 219218 74456 219454
rect 74540 219218 74776 219454
rect 74860 219218 75096 219454
rect 74220 218898 74456 219134
rect 74540 218898 74776 219134
rect 74860 218898 75096 219134
rect 516852 219218 517088 219454
rect 517172 219218 517408 219454
rect 517492 219218 517728 219454
rect 516852 218898 517088 219134
rect 517172 218898 517408 219134
rect 517492 218898 517728 219134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 72860 201218 73096 201454
rect 73180 201218 73416 201454
rect 73500 201218 73736 201454
rect 72860 200898 73096 201134
rect 73180 200898 73416 201134
rect 73500 200898 73736 201134
rect 518212 201218 518448 201454
rect 518532 201218 518768 201454
rect 518852 201218 519088 201454
rect 518212 200898 518448 201134
rect 518532 200898 518768 201134
rect 518852 200898 519088 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 74220 183218 74456 183454
rect 74540 183218 74776 183454
rect 74860 183218 75096 183454
rect 74220 182898 74456 183134
rect 74540 182898 74776 183134
rect 74860 182898 75096 183134
rect 516852 183218 517088 183454
rect 517172 183218 517408 183454
rect 517492 183218 517728 183454
rect 516852 182898 517088 183134
rect 517172 182898 517408 183134
rect 517492 182898 517728 183134
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 72860 165218 73096 165454
rect 73180 165218 73416 165454
rect 73500 165218 73736 165454
rect 72860 164898 73096 165134
rect 73180 164898 73416 165134
rect 73500 164898 73736 165134
rect 518212 165218 518448 165454
rect 518532 165218 518768 165454
rect 518852 165218 519088 165454
rect 518212 164898 518448 165134
rect 518532 164898 518768 165134
rect 518852 164898 519088 165134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 74220 147218 74456 147454
rect 74540 147218 74776 147454
rect 74860 147218 75096 147454
rect 74220 146898 74456 147134
rect 74540 146898 74776 147134
rect 74860 146898 75096 147134
rect 516852 147218 517088 147454
rect 517172 147218 517408 147454
rect 517492 147218 517728 147454
rect 516852 146898 517088 147134
rect 517172 146898 517408 147134
rect 517492 146898 517728 147134
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 72860 129218 73096 129454
rect 73180 129218 73416 129454
rect 73500 129218 73736 129454
rect 72860 128898 73096 129134
rect 73180 128898 73416 129134
rect 73500 128898 73736 129134
rect 518212 129218 518448 129454
rect 518532 129218 518768 129454
rect 518852 129218 519088 129454
rect 518212 128898 518448 129134
rect 518532 128898 518768 129134
rect 518852 128898 519088 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 74220 111218 74456 111454
rect 74540 111218 74776 111454
rect 74860 111218 75096 111454
rect 74220 110898 74456 111134
rect 74540 110898 74776 111134
rect 74860 110898 75096 111134
rect 516852 111218 517088 111454
rect 517172 111218 517408 111454
rect 517492 111218 517728 111454
rect 516852 110898 517088 111134
rect 517172 110898 517408 111134
rect 517492 110898 517728 111134
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 72860 93218 73096 93454
rect 73180 93218 73416 93454
rect 73500 93218 73736 93454
rect 72860 92898 73096 93134
rect 73180 92898 73416 93134
rect 73500 92898 73736 93134
rect 518212 93218 518448 93454
rect 518532 93218 518768 93454
rect 518852 93218 519088 93454
rect 518212 92898 518448 93134
rect 518532 92898 518768 93134
rect 518852 92898 519088 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 74220 75218 74456 75454
rect 74540 75218 74776 75454
rect 74860 75218 75096 75454
rect 74220 74898 74456 75134
rect 74540 74898 74776 75134
rect 74860 74898 75096 75134
rect 516852 75218 517088 75454
rect 517172 75218 517408 75454
rect 517492 75218 517728 75454
rect 516852 74898 517088 75134
rect 517172 74898 517408 75134
rect 517492 74898 517728 75134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 72860 633454
rect 73096 633218 73180 633454
rect 73416 633218 73500 633454
rect 73736 633218 518212 633454
rect 518448 633218 518532 633454
rect 518768 633218 518852 633454
rect 519088 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 72860 633134
rect 73096 632898 73180 633134
rect 73416 632898 73500 633134
rect 73736 632898 518212 633134
rect 518448 632898 518532 633134
rect 518768 632898 518852 633134
rect 519088 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 74220 615454
rect 74456 615218 74540 615454
rect 74776 615218 74860 615454
rect 75096 615218 516852 615454
rect 517088 615218 517172 615454
rect 517408 615218 517492 615454
rect 517728 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 74220 615134
rect 74456 614898 74540 615134
rect 74776 614898 74860 615134
rect 75096 614898 516852 615134
rect 517088 614898 517172 615134
rect 517408 614898 517492 615134
rect 517728 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 72860 597454
rect 73096 597218 73180 597454
rect 73416 597218 73500 597454
rect 73736 597218 518212 597454
rect 518448 597218 518532 597454
rect 518768 597218 518852 597454
rect 519088 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 72860 597134
rect 73096 596898 73180 597134
rect 73416 596898 73500 597134
rect 73736 596898 518212 597134
rect 518448 596898 518532 597134
rect 518768 596898 518852 597134
rect 519088 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 74220 579454
rect 74456 579218 74540 579454
rect 74776 579218 74860 579454
rect 75096 579218 516852 579454
rect 517088 579218 517172 579454
rect 517408 579218 517492 579454
rect 517728 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 74220 579134
rect 74456 578898 74540 579134
rect 74776 578898 74860 579134
rect 75096 578898 516852 579134
rect 517088 578898 517172 579134
rect 517408 578898 517492 579134
rect 517728 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 72860 561454
rect 73096 561218 73180 561454
rect 73416 561218 73500 561454
rect 73736 561218 518212 561454
rect 518448 561218 518532 561454
rect 518768 561218 518852 561454
rect 519088 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 72860 561134
rect 73096 560898 73180 561134
rect 73416 560898 73500 561134
rect 73736 560898 518212 561134
rect 518448 560898 518532 561134
rect 518768 560898 518852 561134
rect 519088 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 74220 543454
rect 74456 543218 74540 543454
rect 74776 543218 74860 543454
rect 75096 543218 516852 543454
rect 517088 543218 517172 543454
rect 517408 543218 517492 543454
rect 517728 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 74220 543134
rect 74456 542898 74540 543134
rect 74776 542898 74860 543134
rect 75096 542898 516852 543134
rect 517088 542898 517172 543134
rect 517408 542898 517492 543134
rect 517728 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 72860 525454
rect 73096 525218 73180 525454
rect 73416 525218 73500 525454
rect 73736 525218 518212 525454
rect 518448 525218 518532 525454
rect 518768 525218 518852 525454
rect 519088 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 72860 525134
rect 73096 524898 73180 525134
rect 73416 524898 73500 525134
rect 73736 524898 518212 525134
rect 518448 524898 518532 525134
rect 518768 524898 518852 525134
rect 519088 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 74220 507454
rect 74456 507218 74540 507454
rect 74776 507218 74860 507454
rect 75096 507218 516852 507454
rect 517088 507218 517172 507454
rect 517408 507218 517492 507454
rect 517728 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 74220 507134
rect 74456 506898 74540 507134
rect 74776 506898 74860 507134
rect 75096 506898 516852 507134
rect 517088 506898 517172 507134
rect 517408 506898 517492 507134
rect 517728 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 72860 489454
rect 73096 489218 73180 489454
rect 73416 489218 73500 489454
rect 73736 489218 518212 489454
rect 518448 489218 518532 489454
rect 518768 489218 518852 489454
rect 519088 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 72860 489134
rect 73096 488898 73180 489134
rect 73416 488898 73500 489134
rect 73736 488898 518212 489134
rect 518448 488898 518532 489134
rect 518768 488898 518852 489134
rect 519088 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 74220 471454
rect 74456 471218 74540 471454
rect 74776 471218 74860 471454
rect 75096 471218 516852 471454
rect 517088 471218 517172 471454
rect 517408 471218 517492 471454
rect 517728 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 74220 471134
rect 74456 470898 74540 471134
rect 74776 470898 74860 471134
rect 75096 470898 516852 471134
rect 517088 470898 517172 471134
rect 517408 470898 517492 471134
rect 517728 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 72860 453454
rect 73096 453218 73180 453454
rect 73416 453218 73500 453454
rect 73736 453218 518212 453454
rect 518448 453218 518532 453454
rect 518768 453218 518852 453454
rect 519088 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 72860 453134
rect 73096 452898 73180 453134
rect 73416 452898 73500 453134
rect 73736 452898 518212 453134
rect 518448 452898 518532 453134
rect 518768 452898 518852 453134
rect 519088 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 74220 435454
rect 74456 435218 74540 435454
rect 74776 435218 74860 435454
rect 75096 435218 516852 435454
rect 517088 435218 517172 435454
rect 517408 435218 517492 435454
rect 517728 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 74220 435134
rect 74456 434898 74540 435134
rect 74776 434898 74860 435134
rect 75096 434898 516852 435134
rect 517088 434898 517172 435134
rect 517408 434898 517492 435134
rect 517728 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 72860 417454
rect 73096 417218 73180 417454
rect 73416 417218 73500 417454
rect 73736 417218 518212 417454
rect 518448 417218 518532 417454
rect 518768 417218 518852 417454
rect 519088 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 72860 417134
rect 73096 416898 73180 417134
rect 73416 416898 73500 417134
rect 73736 416898 518212 417134
rect 518448 416898 518532 417134
rect 518768 416898 518852 417134
rect 519088 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 74220 399454
rect 74456 399218 74540 399454
rect 74776 399218 74860 399454
rect 75096 399218 516852 399454
rect 517088 399218 517172 399454
rect 517408 399218 517492 399454
rect 517728 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 74220 399134
rect 74456 398898 74540 399134
rect 74776 398898 74860 399134
rect 75096 398898 516852 399134
rect 517088 398898 517172 399134
rect 517408 398898 517492 399134
rect 517728 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 72860 381454
rect 73096 381218 73180 381454
rect 73416 381218 73500 381454
rect 73736 381218 518212 381454
rect 518448 381218 518532 381454
rect 518768 381218 518852 381454
rect 519088 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 72860 381134
rect 73096 380898 73180 381134
rect 73416 380898 73500 381134
rect 73736 380898 518212 381134
rect 518448 380898 518532 381134
rect 518768 380898 518852 381134
rect 519088 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74220 363454
rect 74456 363218 74540 363454
rect 74776 363218 74860 363454
rect 75096 363218 516852 363454
rect 517088 363218 517172 363454
rect 517408 363218 517492 363454
rect 517728 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74220 363134
rect 74456 362898 74540 363134
rect 74776 362898 74860 363134
rect 75096 362898 516852 363134
rect 517088 362898 517172 363134
rect 517408 362898 517492 363134
rect 517728 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 72860 345454
rect 73096 345218 73180 345454
rect 73416 345218 73500 345454
rect 73736 345218 518212 345454
rect 518448 345218 518532 345454
rect 518768 345218 518852 345454
rect 519088 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 72860 345134
rect 73096 344898 73180 345134
rect 73416 344898 73500 345134
rect 73736 344898 518212 345134
rect 518448 344898 518532 345134
rect 518768 344898 518852 345134
rect 519088 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 74220 327454
rect 74456 327218 74540 327454
rect 74776 327218 74860 327454
rect 75096 327218 516852 327454
rect 517088 327218 517172 327454
rect 517408 327218 517492 327454
rect 517728 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 74220 327134
rect 74456 326898 74540 327134
rect 74776 326898 74860 327134
rect 75096 326898 516852 327134
rect 517088 326898 517172 327134
rect 517408 326898 517492 327134
rect 517728 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 72860 309454
rect 73096 309218 73180 309454
rect 73416 309218 73500 309454
rect 73736 309218 518212 309454
rect 518448 309218 518532 309454
rect 518768 309218 518852 309454
rect 519088 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 72860 309134
rect 73096 308898 73180 309134
rect 73416 308898 73500 309134
rect 73736 308898 518212 309134
rect 518448 308898 518532 309134
rect 518768 308898 518852 309134
rect 519088 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 74220 291454
rect 74456 291218 74540 291454
rect 74776 291218 74860 291454
rect 75096 291218 516852 291454
rect 517088 291218 517172 291454
rect 517408 291218 517492 291454
rect 517728 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 74220 291134
rect 74456 290898 74540 291134
rect 74776 290898 74860 291134
rect 75096 290898 516852 291134
rect 517088 290898 517172 291134
rect 517408 290898 517492 291134
rect 517728 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 72860 273454
rect 73096 273218 73180 273454
rect 73416 273218 73500 273454
rect 73736 273218 518212 273454
rect 518448 273218 518532 273454
rect 518768 273218 518852 273454
rect 519088 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 72860 273134
rect 73096 272898 73180 273134
rect 73416 272898 73500 273134
rect 73736 272898 518212 273134
rect 518448 272898 518532 273134
rect 518768 272898 518852 273134
rect 519088 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74220 255454
rect 74456 255218 74540 255454
rect 74776 255218 74860 255454
rect 75096 255218 516852 255454
rect 517088 255218 517172 255454
rect 517408 255218 517492 255454
rect 517728 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74220 255134
rect 74456 254898 74540 255134
rect 74776 254898 74860 255134
rect 75096 254898 516852 255134
rect 517088 254898 517172 255134
rect 517408 254898 517492 255134
rect 517728 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 72860 237454
rect 73096 237218 73180 237454
rect 73416 237218 73500 237454
rect 73736 237218 518212 237454
rect 518448 237218 518532 237454
rect 518768 237218 518852 237454
rect 519088 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 72860 237134
rect 73096 236898 73180 237134
rect 73416 236898 73500 237134
rect 73736 236898 518212 237134
rect 518448 236898 518532 237134
rect 518768 236898 518852 237134
rect 519088 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 74220 219454
rect 74456 219218 74540 219454
rect 74776 219218 74860 219454
rect 75096 219218 516852 219454
rect 517088 219218 517172 219454
rect 517408 219218 517492 219454
rect 517728 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 74220 219134
rect 74456 218898 74540 219134
rect 74776 218898 74860 219134
rect 75096 218898 516852 219134
rect 517088 218898 517172 219134
rect 517408 218898 517492 219134
rect 517728 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 72860 201454
rect 73096 201218 73180 201454
rect 73416 201218 73500 201454
rect 73736 201218 518212 201454
rect 518448 201218 518532 201454
rect 518768 201218 518852 201454
rect 519088 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 72860 201134
rect 73096 200898 73180 201134
rect 73416 200898 73500 201134
rect 73736 200898 518212 201134
rect 518448 200898 518532 201134
rect 518768 200898 518852 201134
rect 519088 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 74220 183454
rect 74456 183218 74540 183454
rect 74776 183218 74860 183454
rect 75096 183218 516852 183454
rect 517088 183218 517172 183454
rect 517408 183218 517492 183454
rect 517728 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 74220 183134
rect 74456 182898 74540 183134
rect 74776 182898 74860 183134
rect 75096 182898 516852 183134
rect 517088 182898 517172 183134
rect 517408 182898 517492 183134
rect 517728 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 72860 165454
rect 73096 165218 73180 165454
rect 73416 165218 73500 165454
rect 73736 165218 518212 165454
rect 518448 165218 518532 165454
rect 518768 165218 518852 165454
rect 519088 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 72860 165134
rect 73096 164898 73180 165134
rect 73416 164898 73500 165134
rect 73736 164898 518212 165134
rect 518448 164898 518532 165134
rect 518768 164898 518852 165134
rect 519088 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 74220 147454
rect 74456 147218 74540 147454
rect 74776 147218 74860 147454
rect 75096 147218 516852 147454
rect 517088 147218 517172 147454
rect 517408 147218 517492 147454
rect 517728 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 74220 147134
rect 74456 146898 74540 147134
rect 74776 146898 74860 147134
rect 75096 146898 516852 147134
rect 517088 146898 517172 147134
rect 517408 146898 517492 147134
rect 517728 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 72860 129454
rect 73096 129218 73180 129454
rect 73416 129218 73500 129454
rect 73736 129218 518212 129454
rect 518448 129218 518532 129454
rect 518768 129218 518852 129454
rect 519088 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 72860 129134
rect 73096 128898 73180 129134
rect 73416 128898 73500 129134
rect 73736 128898 518212 129134
rect 518448 128898 518532 129134
rect 518768 128898 518852 129134
rect 519088 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 74220 111454
rect 74456 111218 74540 111454
rect 74776 111218 74860 111454
rect 75096 111218 516852 111454
rect 517088 111218 517172 111454
rect 517408 111218 517492 111454
rect 517728 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 74220 111134
rect 74456 110898 74540 111134
rect 74776 110898 74860 111134
rect 75096 110898 516852 111134
rect 517088 110898 517172 111134
rect 517408 110898 517492 111134
rect 517728 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 72860 93454
rect 73096 93218 73180 93454
rect 73416 93218 73500 93454
rect 73736 93218 518212 93454
rect 518448 93218 518532 93454
rect 518768 93218 518852 93454
rect 519088 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 72860 93134
rect 73096 92898 73180 93134
rect 73416 92898 73500 93134
rect 73736 92898 518212 93134
rect 518448 92898 518532 93134
rect 518768 92898 518852 93134
rect 519088 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 74220 75454
rect 74456 75218 74540 75454
rect 74776 75218 74860 75454
rect 75096 75218 516852 75454
rect 517088 75218 517172 75454
rect 517408 75218 517492 75454
rect 517728 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 74220 75134
rect 74456 74898 74540 75134
rect 74776 74898 74860 75134
rect 75096 74898 516852 75134
rect 517088 74898 517172 75134
rect 517408 74898 517492 75134
rect 517728 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Ibtida_top_dffram_cv  mprj
timestamp 1635531245
transform 1 0 72000 0 1 60000
box 0 0 447948 592008
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 654008 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 654008 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 654008 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 654008 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 654008 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 654008 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 654008 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 654008 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 654008 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 654008 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 654008 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 654008 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 654008 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 654008 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 654008 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 654008 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 654008 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 654008 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 654008 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 654008 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 654008 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 654008 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 654008 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 654008 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 654008 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 654008 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 654008 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 654008 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 654008 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 654008 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 654008 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 654008 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 654008 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 654008 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 654008 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 654008 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 654008 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 654008 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 654008 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 654008 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 654008 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 654008 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 654008 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 654008 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 654008 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 654008 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 654008 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 654008 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 654008 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 654008 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 654008 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 654008 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 654008 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 654008 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 654008 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 654008 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 654008 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 654008 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 654008 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 654008 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 654008 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 654008 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 654008 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 654008 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 654008 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 654008 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 654008 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 654008 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 654008 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 654008 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 654008 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 654008 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 654008 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 654008 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 654008 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 654008 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 654008 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 654008 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 654008 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 654008 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 654008 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 654008 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 654008 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 654008 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 654008 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 654008 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 654008 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 654008 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 654008 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 654008 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 654008 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 654008 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 654008 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 654008 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 654008 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 654008 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 654008 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 654008 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 654008 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 654008 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
