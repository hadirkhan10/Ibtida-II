##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Oct 29 16:53:51 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Ibtida_top_dffram_cv
  CLASS BLOCK ;
  SIZE 2239.740000 BY 2960.040000 ;
  FOREIGN Ibtida_top_dffram_cv 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760000 0.000000 4.900000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300000 0.000000 4.440000 0.490000 ;
    END
  END wb_rst_i
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.160000 0.000000 1058.300000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.560000 0.000000 1053.700000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.960000 0.000000 1049.100000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.820000 0.000000 1044.960000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.220000 0.000000 1040.360000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.620000 0.000000 1035.760000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.020000 0.000000 1031.160000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.420000 0.000000 1026.560000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.820000 0.000000 1021.960000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.220000 0.000000 1017.360000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.620000 0.000000 1012.760000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.020000 0.000000 1008.160000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.880000 0.000000 1004.020000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.280000 0.000000 999.420000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.680000 0.000000 994.820000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.080000 0.000000 990.220000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.480000 0.000000 985.620000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.880000 0.000000 981.020000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.280000 0.000000 976.420000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.680000 0.000000 971.820000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.540000 0.000000 967.680000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.940000 0.000000 963.080000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.340000 0.000000 958.480000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.740000 0.000000 953.880000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.140000 0.000000 949.280000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.540000 0.000000 944.680000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.940000 0.000000 940.080000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.340000 0.000000 935.480000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.200000 0.000000 931.340000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.600000 0.000000 926.740000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.000000 0.000000 922.140000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.400000 0.000000 917.540000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.800000 0.000000 912.940000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.200000 0.000000 908.340000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.600000 0.000000 903.740000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.000000 0.000000 899.140000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.860000 0.000000 895.000000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.260000 0.000000 890.400000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.660000 0.000000 885.800000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.060000 0.000000 881.200000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.460000 0.000000 876.600000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.860000 0.000000 872.000000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.260000 0.000000 867.400000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.660000 0.000000 862.800000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.520000 0.000000 858.660000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.920000 0.000000 854.060000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.320000 0.000000 849.460000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.720000 0.000000 844.860000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.120000 0.000000 840.260000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.520000 0.000000 835.660000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.920000 0.000000 831.060000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.320000 0.000000 826.460000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.180000 0.000000 822.320000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.580000 0.000000 817.720000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.980000 0.000000 813.120000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.380000 0.000000 808.520000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.780000 0.000000 803.920000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.180000 0.000000 799.320000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.580000 0.000000 794.720000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.980000 0.000000 790.120000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.840000 0.000000 785.980000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.240000 0.000000 781.380000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.640000 0.000000 776.780000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.040000 0.000000 772.180000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.440000 0.000000 767.580000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.840000 0.000000 762.980000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.240000 0.000000 758.380000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.640000 0.000000 753.780000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.500000 0.000000 749.640000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.900000 0.000000 745.040000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.300000 0.000000 740.440000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.700000 0.000000 735.840000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.100000 0.000000 731.240000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.500000 0.000000 726.640000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.900000 0.000000 722.040000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.300000 0.000000 717.440000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.160000 0.000000 713.300000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.560000 0.000000 708.700000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.960000 0.000000 704.100000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.360000 0.000000 699.500000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.760000 0.000000 694.900000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.160000 0.000000 690.300000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.560000 0.000000 685.700000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.960000 0.000000 681.100000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.820000 0.000000 676.960000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.220000 0.000000 672.360000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.620000 0.000000 667.760000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.020000 0.000000 663.160000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.420000 0.000000 658.560000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.820000 0.000000 653.960000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.220000 0.000000 649.360000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.620000 0.000000 644.760000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.480000 0.000000 640.620000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.880000 0.000000 636.020000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.280000 0.000000 631.420000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.680000 0.000000 626.820000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.080000 0.000000 622.220000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.480000 0.000000 617.620000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.880000 0.000000 613.020000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.280000 0.000000 608.420000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.140000 0.000000 604.280000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.540000 0.000000 599.680000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.940000 0.000000 595.080000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.340000 0.000000 590.480000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.740000 0.000000 585.880000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.140000 0.000000 581.280000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.540000 0.000000 576.680000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.940000 0.000000 572.080000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.800000 0.000000 567.940000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.200000 0.000000 563.340000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.600000 0.000000 558.740000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.000000 0.000000 554.140000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.400000 0.000000 549.540000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.800000 0.000000 544.940000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.200000 0.000000 540.340000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.600000 0.000000 535.740000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.460000 0.000000 531.600000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.860000 0.000000 527.000000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.260000 0.000000 522.400000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.660000 0.000000 517.800000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.060000 0.000000 513.200000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.460000 0.000000 508.600000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.860000 0.000000 504.000000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.260000 0.000000 499.400000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.660000 0.000000 494.800000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.520000 0.000000 490.660000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.920000 0.000000 486.060000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.320000 0.000000 481.460000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.600000 0.000000 1639.740000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.000000 0.000000 1635.140000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.860000 0.000000 1631.000000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.260000 0.000000 1626.400000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.660000 0.000000 1621.800000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.060000 0.000000 1617.200000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.460000 0.000000 1612.600000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.860000 0.000000 1608.000000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.260000 0.000000 1603.400000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.660000 0.000000 1598.800000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.520000 0.000000 1594.660000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.920000 0.000000 1590.060000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.320000 0.000000 1585.460000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.720000 0.000000 1580.860000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.120000 0.000000 1576.260000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.520000 0.000000 1571.660000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.920000 0.000000 1567.060000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.320000 0.000000 1562.460000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.180000 0.000000 1558.320000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.580000 0.000000 1553.720000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.980000 0.000000 1549.120000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.380000 0.000000 1544.520000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.780000 0.000000 1539.920000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.180000 0.000000 1535.320000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.580000 0.000000 1530.720000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.980000 0.000000 1526.120000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.380000 0.000000 1521.520000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.240000 0.000000 1517.380000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.640000 0.000000 1512.780000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.040000 0.000000 1508.180000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.440000 0.000000 1503.580000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.840000 0.000000 1498.980000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.240000 0.000000 1494.380000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.640000 0.000000 1489.780000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.040000 0.000000 1485.180000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.900000 0.000000 1481.040000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.300000 0.000000 1476.440000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.700000 0.000000 1471.840000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.100000 0.000000 1467.240000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.500000 0.000000 1462.640000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.900000 0.000000 1458.040000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.300000 0.000000 1453.440000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.700000 0.000000 1448.840000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.560000 0.000000 1444.700000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.960000 0.000000 1440.100000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.360000 0.000000 1435.500000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.760000 0.000000 1430.900000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.160000 0.000000 1426.300000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.560000 0.000000 1421.700000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.960000 0.000000 1417.100000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.360000 0.000000 1412.500000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.220000 0.000000 1408.360000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.620000 0.000000 1403.760000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.020000 0.000000 1399.160000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.420000 0.000000 1394.560000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.820000 0.000000 1389.960000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.220000 0.000000 1385.360000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.620000 0.000000 1380.760000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.020000 0.000000 1376.160000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.880000 0.000000 1372.020000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.280000 0.000000 1367.420000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.680000 0.000000 1362.820000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.080000 0.000000 1358.220000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.480000 0.000000 1353.620000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.880000 0.000000 1349.020000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.280000 0.000000 1344.420000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.680000 0.000000 1339.820000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.540000 0.000000 1335.680000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.940000 0.000000 1331.080000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.340000 0.000000 1326.480000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.740000 0.000000 1321.880000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.140000 0.000000 1317.280000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.540000 0.000000 1312.680000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.940000 0.000000 1308.080000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.340000 0.000000 1303.480000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.200000 0.000000 1299.340000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.600000 0.000000 1294.740000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.000000 0.000000 1290.140000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.400000 0.000000 1285.540000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.800000 0.000000 1280.940000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.200000 0.000000 1276.340000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.600000 0.000000 1271.740000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.000000 0.000000 1267.140000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.860000 0.000000 1263.000000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.260000 0.000000 1258.400000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.660000 0.000000 1253.800000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.060000 0.000000 1249.200000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.460000 0.000000 1244.600000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.860000 0.000000 1240.000000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.260000 0.000000 1235.400000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.660000 0.000000 1230.800000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.520000 0.000000 1226.660000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.920000 0.000000 1222.060000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.320000 0.000000 1217.460000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.720000 0.000000 1212.860000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.120000 0.000000 1208.260000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.520000 0.000000 1203.660000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.920000 0.000000 1199.060000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.320000 0.000000 1194.460000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.180000 0.000000 1190.320000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.580000 0.000000 1185.720000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.980000 0.000000 1181.120000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.380000 0.000000 1176.520000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.780000 0.000000 1171.920000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.180000 0.000000 1167.320000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.580000 0.000000 1162.720000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.980000 0.000000 1158.120000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.840000 0.000000 1153.980000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.240000 0.000000 1149.380000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.640000 0.000000 1144.780000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.040000 0.000000 1140.180000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.440000 0.000000 1135.580000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.840000 0.000000 1130.980000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.240000 0.000000 1126.380000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.640000 0.000000 1121.780000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.500000 0.000000 1117.640000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.900000 0.000000 1113.040000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.300000 0.000000 1108.440000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.700000 0.000000 1103.840000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.100000 0.000000 1099.240000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.500000 0.000000 1094.640000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.900000 0.000000 1090.040000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.300000 0.000000 1085.440000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.160000 0.000000 1081.300000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.560000 0.000000 1076.700000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.960000 0.000000 1072.100000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.360000 0.000000 1067.500000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.760000 0.000000 1062.900000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.040000 0.000000 2221.180000 0.490000 ;
    END
  END la_oen[127]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.900000 0.000000 2217.040000 0.490000 ;
    END
  END la_oen[126]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.300000 0.000000 2212.440000 0.490000 ;
    END
  END la_oen[125]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.700000 0.000000 2207.840000 0.490000 ;
    END
  END la_oen[124]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.100000 0.000000 2203.240000 0.490000 ;
    END
  END la_oen[123]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.500000 0.000000 2198.640000 0.490000 ;
    END
  END la_oen[122]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.900000 0.000000 2194.040000 0.490000 ;
    END
  END la_oen[121]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.300000 0.000000 2189.440000 0.490000 ;
    END
  END la_oen[120]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.700000 0.000000 2184.840000 0.490000 ;
    END
  END la_oen[119]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.560000 0.000000 2180.700000 0.490000 ;
    END
  END la_oen[118]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.960000 0.000000 2176.100000 0.490000 ;
    END
  END la_oen[117]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.360000 0.000000 2171.500000 0.490000 ;
    END
  END la_oen[116]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.760000 0.000000 2166.900000 0.490000 ;
    END
  END la_oen[115]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.160000 0.000000 2162.300000 0.490000 ;
    END
  END la_oen[114]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.560000 0.000000 2157.700000 0.490000 ;
    END
  END la_oen[113]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.960000 0.000000 2153.100000 0.490000 ;
    END
  END la_oen[112]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.360000 0.000000 2148.500000 0.490000 ;
    END
  END la_oen[111]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.220000 0.000000 2144.360000 0.490000 ;
    END
  END la_oen[110]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.620000 0.000000 2139.760000 0.490000 ;
    END
  END la_oen[109]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.020000 0.000000 2135.160000 0.490000 ;
    END
  END la_oen[108]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.420000 0.000000 2130.560000 0.490000 ;
    END
  END la_oen[107]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.820000 0.000000 2125.960000 0.490000 ;
    END
  END la_oen[106]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.220000 0.000000 2121.360000 0.490000 ;
    END
  END la_oen[105]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.620000 0.000000 2116.760000 0.490000 ;
    END
  END la_oen[104]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.020000 0.000000 2112.160000 0.490000 ;
    END
  END la_oen[103]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.880000 0.000000 2108.020000 0.490000 ;
    END
  END la_oen[102]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.280000 0.000000 2103.420000 0.490000 ;
    END
  END la_oen[101]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.680000 0.000000 2098.820000 0.490000 ;
    END
  END la_oen[100]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.080000 0.000000 2094.220000 0.490000 ;
    END
  END la_oen[99]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.480000 0.000000 2089.620000 0.490000 ;
    END
  END la_oen[98]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.880000 0.000000 2085.020000 0.490000 ;
    END
  END la_oen[97]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.280000 0.000000 2080.420000 0.490000 ;
    END
  END la_oen[96]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.680000 0.000000 2075.820000 0.490000 ;
    END
  END la_oen[95]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.540000 0.000000 2071.680000 0.490000 ;
    END
  END la_oen[94]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.940000 0.000000 2067.080000 0.490000 ;
    END
  END la_oen[93]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.340000 0.000000 2062.480000 0.490000 ;
    END
  END la_oen[92]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.740000 0.000000 2057.880000 0.490000 ;
    END
  END la_oen[91]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.140000 0.000000 2053.280000 0.490000 ;
    END
  END la_oen[90]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.540000 0.000000 2048.680000 0.490000 ;
    END
  END la_oen[89]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.940000 0.000000 2044.080000 0.490000 ;
    END
  END la_oen[88]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.340000 0.000000 2039.480000 0.490000 ;
    END
  END la_oen[87]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.740000 0.000000 2034.880000 0.490000 ;
    END
  END la_oen[86]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.600000 0.000000 2030.740000 0.490000 ;
    END
  END la_oen[85]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.000000 0.000000 2026.140000 0.490000 ;
    END
  END la_oen[84]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.400000 0.000000 2021.540000 0.490000 ;
    END
  END la_oen[83]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.800000 0.000000 2016.940000 0.490000 ;
    END
  END la_oen[82]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.200000 0.000000 2012.340000 0.490000 ;
    END
  END la_oen[81]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.600000 0.000000 2007.740000 0.490000 ;
    END
  END la_oen[80]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.000000 0.000000 2003.140000 0.490000 ;
    END
  END la_oen[79]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.400000 0.000000 1998.540000 0.490000 ;
    END
  END la_oen[78]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.260000 0.000000 1994.400000 0.490000 ;
    END
  END la_oen[77]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.660000 0.000000 1989.800000 0.490000 ;
    END
  END la_oen[76]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.060000 0.000000 1985.200000 0.490000 ;
    END
  END la_oen[75]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.460000 0.000000 1980.600000 0.490000 ;
    END
  END la_oen[74]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.860000 0.000000 1976.000000 0.490000 ;
    END
  END la_oen[73]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.260000 0.000000 1971.400000 0.490000 ;
    END
  END la_oen[72]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.660000 0.000000 1966.800000 0.490000 ;
    END
  END la_oen[71]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.060000 0.000000 1962.200000 0.490000 ;
    END
  END la_oen[70]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.920000 0.000000 1958.060000 0.490000 ;
    END
  END la_oen[69]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.320000 0.000000 1953.460000 0.490000 ;
    END
  END la_oen[68]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.720000 0.000000 1948.860000 0.490000 ;
    END
  END la_oen[67]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.120000 0.000000 1944.260000 0.490000 ;
    END
  END la_oen[66]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.520000 0.000000 1939.660000 0.490000 ;
    END
  END la_oen[65]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.920000 0.000000 1935.060000 0.490000 ;
    END
  END la_oen[64]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.320000 0.000000 1930.460000 0.490000 ;
    END
  END la_oen[63]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.720000 0.000000 1925.860000 0.490000 ;
    END
  END la_oen[62]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.580000 0.000000 1921.720000 0.490000 ;
    END
  END la_oen[61]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.980000 0.000000 1917.120000 0.490000 ;
    END
  END la_oen[60]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.380000 0.000000 1912.520000 0.490000 ;
    END
  END la_oen[59]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.780000 0.000000 1907.920000 0.490000 ;
    END
  END la_oen[58]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.180000 0.000000 1903.320000 0.490000 ;
    END
  END la_oen[57]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.580000 0.000000 1898.720000 0.490000 ;
    END
  END la_oen[56]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.980000 0.000000 1894.120000 0.490000 ;
    END
  END la_oen[55]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.380000 0.000000 1889.520000 0.490000 ;
    END
  END la_oen[54]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.240000 0.000000 1885.380000 0.490000 ;
    END
  END la_oen[53]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.640000 0.000000 1880.780000 0.490000 ;
    END
  END la_oen[52]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.040000 0.000000 1876.180000 0.490000 ;
    END
  END la_oen[51]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.440000 0.000000 1871.580000 0.490000 ;
    END
  END la_oen[50]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.840000 0.000000 1866.980000 0.490000 ;
    END
  END la_oen[49]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.240000 0.000000 1862.380000 0.490000 ;
    END
  END la_oen[48]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.640000 0.000000 1857.780000 0.490000 ;
    END
  END la_oen[47]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.040000 0.000000 1853.180000 0.490000 ;
    END
  END la_oen[46]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.900000 0.000000 1849.040000 0.490000 ;
    END
  END la_oen[45]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.300000 0.000000 1844.440000 0.490000 ;
    END
  END la_oen[44]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.700000 0.000000 1839.840000 0.490000 ;
    END
  END la_oen[43]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.100000 0.000000 1835.240000 0.490000 ;
    END
  END la_oen[42]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.500000 0.000000 1830.640000 0.490000 ;
    END
  END la_oen[41]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.900000 0.000000 1826.040000 0.490000 ;
    END
  END la_oen[40]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.300000 0.000000 1821.440000 0.490000 ;
    END
  END la_oen[39]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.700000 0.000000 1816.840000 0.490000 ;
    END
  END la_oen[38]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.560000 0.000000 1812.700000 0.490000 ;
    END
  END la_oen[37]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.960000 0.000000 1808.100000 0.490000 ;
    END
  END la_oen[36]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.360000 0.000000 1803.500000 0.490000 ;
    END
  END la_oen[35]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.760000 0.000000 1798.900000 0.490000 ;
    END
  END la_oen[34]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.160000 0.000000 1794.300000 0.490000 ;
    END
  END la_oen[33]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.560000 0.000000 1789.700000 0.490000 ;
    END
  END la_oen[32]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.960000 0.000000 1785.100000 0.490000 ;
    END
  END la_oen[31]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.360000 0.000000 1780.500000 0.490000 ;
    END
  END la_oen[30]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.220000 0.000000 1776.360000 0.490000 ;
    END
  END la_oen[29]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.620000 0.000000 1771.760000 0.490000 ;
    END
  END la_oen[28]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.020000 0.000000 1767.160000 0.490000 ;
    END
  END la_oen[27]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.420000 0.000000 1762.560000 0.490000 ;
    END
  END la_oen[26]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.820000 0.000000 1757.960000 0.490000 ;
    END
  END la_oen[25]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1753.220000 0.000000 1753.360000 0.490000 ;
    END
  END la_oen[24]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.620000 0.000000 1748.760000 0.490000 ;
    END
  END la_oen[23]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.020000 0.000000 1744.160000 0.490000 ;
    END
  END la_oen[22]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.880000 0.000000 1740.020000 0.490000 ;
    END
  END la_oen[21]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.280000 0.000000 1735.420000 0.490000 ;
    END
  END la_oen[20]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.680000 0.000000 1730.820000 0.490000 ;
    END
  END la_oen[19]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.080000 0.000000 1726.220000 0.490000 ;
    END
  END la_oen[18]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.480000 0.000000 1721.620000 0.490000 ;
    END
  END la_oen[17]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.880000 0.000000 1717.020000 0.490000 ;
    END
  END la_oen[16]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.280000 0.000000 1712.420000 0.490000 ;
    END
  END la_oen[15]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.680000 0.000000 1707.820000 0.490000 ;
    END
  END la_oen[14]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.540000 0.000000 1703.680000 0.490000 ;
    END
  END la_oen[13]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.940000 0.000000 1699.080000 0.490000 ;
    END
  END la_oen[12]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.340000 0.000000 1694.480000 0.490000 ;
    END
  END la_oen[11]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.740000 0.000000 1689.880000 0.490000 ;
    END
  END la_oen[10]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.140000 0.000000 1685.280000 0.490000 ;
    END
  END la_oen[9]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.540000 0.000000 1680.680000 0.490000 ;
    END
  END la_oen[8]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.940000 0.000000 1676.080000 0.490000 ;
    END
  END la_oen[7]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.340000 0.000000 1671.480000 0.490000 ;
    END
  END la_oen[6]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.200000 0.000000 1667.340000 0.490000 ;
    END
  END la_oen[5]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.600000 0.000000 1662.740000 0.490000 ;
    END
  END la_oen[4]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.000000 0.000000 1658.140000 0.490000 ;
    END
  END la_oen[3]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.400000 0.000000 1653.540000 0.490000 ;
    END
  END la_oen[2]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.800000 0.000000 1648.940000 0.490000 ;
    END
  END la_oen[1]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.200000 0.000000 1644.340000 0.490000 ;
    END
  END la_oen[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 111.580000 0.800000 111.880000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 279.330000 0.800000 279.630000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 447.080000 0.800000 447.380000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 670.340000 0.800000 670.640000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 893.600000 0.800000 893.900000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1116.860000 0.800000 1117.160000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1340.730000 0.800000 1341.030000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1563.990000 0.800000 1564.290000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1787.250000 0.800000 1787.550000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2010.510000 0.800000 2010.810000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2234.380000 0.800000 2234.680000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2457.640000 0.800000 2457.940000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2680.900000 0.800000 2681.200000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2904.160000 0.800000 2904.460000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040000 2959.550000 128.180000 2960.040000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.260000 2959.550000 384.400000 2960.040000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.020000 2959.550000 640.160000 2960.040000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.240000 2959.550000 896.380000 2960.040000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.000000 2959.550000 1152.140000 2960.040000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.760000 2959.550000 1407.900000 2960.040000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.980000 2959.550000 1664.120000 2960.040000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.740000 2959.550000 1919.880000 2960.040000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.960000 2959.550000 2176.100000 2960.040000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2845.600000 2239.740000 2845.900000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2618.070000 2239.740000 2618.370000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2390.540000 2239.740000 2390.840000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2162.400000 2239.740000 2162.700000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1934.870000 2239.740000 1935.170000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1707.340000 2239.740000 1707.640000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1479.810000 2239.740000 1480.110000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1251.670000 2239.740000 1251.970000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1024.140000 2239.740000 1024.440000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 853.340000 2239.740000 853.640000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 682.540000 2239.740000 682.840000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 511.740000 2239.740000 512.040000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 340.940000 2239.740000 341.240000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 170.140000 2239.740000 170.440000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 4.220000 2239.740000 4.520000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.070000 0.800000 56.370000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 223.820000 0.800000 224.120000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 390.960000 0.800000 391.260000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 614.220000 0.800000 614.520000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 838.090000 0.800000 838.390000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1061.350000 0.800000 1061.650000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1284.610000 0.800000 1284.910000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1507.870000 0.800000 1508.170000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1731.740000 0.800000 1732.040000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1955.000000 0.800000 1955.300000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2178.260000 0.800000 2178.560000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2401.520000 0.800000 2401.820000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2624.780000 0.800000 2625.080000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2848.650000 0.800000 2848.950000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100000 2959.550000 64.240000 2960.040000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.320000 2959.550000 320.460000 2960.040000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.080000 2959.550000 576.220000 2960.040000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.840000 2959.550000 831.980000 2960.040000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.060000 2959.550000 1088.200000 2960.040000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.820000 2959.550000 1343.960000 2960.040000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.040000 2959.550000 1600.180000 2960.040000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.800000 2959.550000 1855.940000 2960.040000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.020000 2959.550000 2112.160000 2960.040000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2902.330000 2239.740000 2902.630000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2674.800000 2239.740000 2675.100000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2447.270000 2239.740000 2447.570000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2219.740000 2239.740000 2220.040000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1991.600000 2239.740000 1991.900000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1764.070000 2239.740000 1764.370000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1536.540000 2239.740000 1536.840000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1309.010000 2239.740000 1309.310000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1080.870000 2239.740000 1081.170000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 910.070000 2239.740000 910.370000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 739.270000 2239.740000 739.570000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 569.080000 2239.740000 569.380000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 398.280000 2239.740000 398.580000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 227.480000 2239.740000 227.780000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 56.680000 2239.740000 56.980000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.440000 0.800000 5.740000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.700000 0.800000 168.000000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 335.450000 0.800000 335.750000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 558.710000 0.800000 559.010000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 781.970000 0.800000 782.270000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1005.230000 0.800000 1005.530000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1229.100000 0.800000 1229.400000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1452.360000 0.800000 1452.660000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1675.620000 0.800000 1675.920000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1898.880000 0.800000 1899.180000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2122.140000 0.800000 2122.440000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2346.010000 0.800000 2346.310000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2569.270000 0.800000 2569.570000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2792.530000 0.800000 2792.830000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.220000 2959.550000 5.360000 2960.040000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.920000 2959.550000 256.060000 2960.040000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.140000 2959.550000 512.280000 2960.040000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.900000 2959.550000 768.040000 2960.040000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.120000 2959.550000 1024.260000 2960.040000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.880000 2959.550000 1280.020000 2960.040000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.100000 2959.550000 1536.240000 2960.040000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.860000 2959.550000 1792.000000 2960.040000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.080000 2959.550000 2048.220000 2960.040000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2954.180000 2239.740000 2954.480000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2732.140000 2239.740000 2732.440000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2504.000000 2239.740000 2504.300000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2276.470000 2239.740000 2276.770000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 2048.940000 2239.740000 2049.240000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1820.800000 2239.740000 1821.100000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1593.270000 2239.740000 1593.570000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1365.740000 2239.740000 1366.040000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 1138.210000 2239.740000 1138.510000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 967.410000 2239.740000 967.710000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 796.610000 2239.740000 796.910000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 625.810000 2239.740000 626.110000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 455.010000 2239.740000 455.310000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 284.210000 2239.740000 284.510000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2238.940000 113.410000 2239.740000 113.710000 ;
    END
  END io_oeb[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2230.750000 4.130000 2235.750000 2955.230000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.990000 4.130000 8.990000 2955.230000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.790000 10.930000 15.790000 2948.430000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.950000 10.930000 2228.950000 2948.430000 ;
    END
  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2239.740000 2960.040000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2239.740000 2960.040000 ;
    LAYER met2 ;
      RECT 2176.240000 2959.410000 2239.740000 2960.040000 ;
      RECT 2112.300000 2959.410000 2175.820000 2960.040000 ;
      RECT 2048.360000 2959.410000 2111.880000 2960.040000 ;
      RECT 1920.020000 2959.410000 2047.940000 2960.040000 ;
      RECT 1856.080000 2959.410000 1919.600000 2960.040000 ;
      RECT 1792.140000 2959.410000 1855.660000 2960.040000 ;
      RECT 1664.260000 2959.410000 1791.720000 2960.040000 ;
      RECT 1600.320000 2959.410000 1663.840000 2960.040000 ;
      RECT 1536.380000 2959.410000 1599.900000 2960.040000 ;
      RECT 1408.040000 2959.410000 1535.960000 2960.040000 ;
      RECT 1344.100000 2959.410000 1407.620000 2960.040000 ;
      RECT 1280.160000 2959.410000 1343.680000 2960.040000 ;
      RECT 1152.280000 2959.410000 1279.740000 2960.040000 ;
      RECT 1088.340000 2959.410000 1151.860000 2960.040000 ;
      RECT 1024.400000 2959.410000 1087.920000 2960.040000 ;
      RECT 896.520000 2959.410000 1023.980000 2960.040000 ;
      RECT 832.120000 2959.410000 896.100000 2960.040000 ;
      RECT 768.180000 2959.410000 831.700000 2960.040000 ;
      RECT 640.300000 2959.410000 767.760000 2960.040000 ;
      RECT 576.360000 2959.410000 639.880000 2960.040000 ;
      RECT 512.420000 2959.410000 575.940000 2960.040000 ;
      RECT 384.540000 2959.410000 512.000000 2960.040000 ;
      RECT 320.600000 2959.410000 384.120000 2960.040000 ;
      RECT 256.200000 2959.410000 320.180000 2960.040000 ;
      RECT 128.320000 2959.410000 255.780000 2960.040000 ;
      RECT 64.380000 2959.410000 127.900000 2960.040000 ;
      RECT 5.500000 2959.410000 63.960000 2960.040000 ;
      RECT 0.000000 2959.410000 5.080000 2960.040000 ;
      RECT 0.000000 0.630000 2239.740000 2959.410000 ;
      RECT 2221.320000 0.000000 2239.740000 0.630000 ;
      RECT 2217.180000 0.000000 2220.900000 0.630000 ;
      RECT 2212.580000 0.000000 2216.760000 0.630000 ;
      RECT 2207.980000 0.000000 2212.160000 0.630000 ;
      RECT 2203.380000 0.000000 2207.560000 0.630000 ;
      RECT 2198.780000 0.000000 2202.960000 0.630000 ;
      RECT 2194.180000 0.000000 2198.360000 0.630000 ;
      RECT 2189.580000 0.000000 2193.760000 0.630000 ;
      RECT 2184.980000 0.000000 2189.160000 0.630000 ;
      RECT 2180.840000 0.000000 2184.560000 0.630000 ;
      RECT 2176.240000 0.000000 2180.420000 0.630000 ;
      RECT 2171.640000 0.000000 2175.820000 0.630000 ;
      RECT 2167.040000 0.000000 2171.220000 0.630000 ;
      RECT 2162.440000 0.000000 2166.620000 0.630000 ;
      RECT 2157.840000 0.000000 2162.020000 0.630000 ;
      RECT 2153.240000 0.000000 2157.420000 0.630000 ;
      RECT 2148.640000 0.000000 2152.820000 0.630000 ;
      RECT 2144.500000 0.000000 2148.220000 0.630000 ;
      RECT 2139.900000 0.000000 2144.080000 0.630000 ;
      RECT 2135.300000 0.000000 2139.480000 0.630000 ;
      RECT 2130.700000 0.000000 2134.880000 0.630000 ;
      RECT 2126.100000 0.000000 2130.280000 0.630000 ;
      RECT 2121.500000 0.000000 2125.680000 0.630000 ;
      RECT 2116.900000 0.000000 2121.080000 0.630000 ;
      RECT 2112.300000 0.000000 2116.480000 0.630000 ;
      RECT 2108.160000 0.000000 2111.880000 0.630000 ;
      RECT 2103.560000 0.000000 2107.740000 0.630000 ;
      RECT 2098.960000 0.000000 2103.140000 0.630000 ;
      RECT 2094.360000 0.000000 2098.540000 0.630000 ;
      RECT 2089.760000 0.000000 2093.940000 0.630000 ;
      RECT 2085.160000 0.000000 2089.340000 0.630000 ;
      RECT 2080.560000 0.000000 2084.740000 0.630000 ;
      RECT 2075.960000 0.000000 2080.140000 0.630000 ;
      RECT 2071.820000 0.000000 2075.540000 0.630000 ;
      RECT 2067.220000 0.000000 2071.400000 0.630000 ;
      RECT 2062.620000 0.000000 2066.800000 0.630000 ;
      RECT 2058.020000 0.000000 2062.200000 0.630000 ;
      RECT 2053.420000 0.000000 2057.600000 0.630000 ;
      RECT 2048.820000 0.000000 2053.000000 0.630000 ;
      RECT 2044.220000 0.000000 2048.400000 0.630000 ;
      RECT 2039.620000 0.000000 2043.800000 0.630000 ;
      RECT 2035.020000 0.000000 2039.200000 0.630000 ;
      RECT 2030.880000 0.000000 2034.600000 0.630000 ;
      RECT 2026.280000 0.000000 2030.460000 0.630000 ;
      RECT 2021.680000 0.000000 2025.860000 0.630000 ;
      RECT 2017.080000 0.000000 2021.260000 0.630000 ;
      RECT 2012.480000 0.000000 2016.660000 0.630000 ;
      RECT 2007.880000 0.000000 2012.060000 0.630000 ;
      RECT 2003.280000 0.000000 2007.460000 0.630000 ;
      RECT 1998.680000 0.000000 2002.860000 0.630000 ;
      RECT 1994.540000 0.000000 1998.260000 0.630000 ;
      RECT 1989.940000 0.000000 1994.120000 0.630000 ;
      RECT 1985.340000 0.000000 1989.520000 0.630000 ;
      RECT 1980.740000 0.000000 1984.920000 0.630000 ;
      RECT 1976.140000 0.000000 1980.320000 0.630000 ;
      RECT 1971.540000 0.000000 1975.720000 0.630000 ;
      RECT 1966.940000 0.000000 1971.120000 0.630000 ;
      RECT 1962.340000 0.000000 1966.520000 0.630000 ;
      RECT 1958.200000 0.000000 1961.920000 0.630000 ;
      RECT 1953.600000 0.000000 1957.780000 0.630000 ;
      RECT 1949.000000 0.000000 1953.180000 0.630000 ;
      RECT 1944.400000 0.000000 1948.580000 0.630000 ;
      RECT 1939.800000 0.000000 1943.980000 0.630000 ;
      RECT 1935.200000 0.000000 1939.380000 0.630000 ;
      RECT 1930.600000 0.000000 1934.780000 0.630000 ;
      RECT 1926.000000 0.000000 1930.180000 0.630000 ;
      RECT 1921.860000 0.000000 1925.580000 0.630000 ;
      RECT 1917.260000 0.000000 1921.440000 0.630000 ;
      RECT 1912.660000 0.000000 1916.840000 0.630000 ;
      RECT 1908.060000 0.000000 1912.240000 0.630000 ;
      RECT 1903.460000 0.000000 1907.640000 0.630000 ;
      RECT 1898.860000 0.000000 1903.040000 0.630000 ;
      RECT 1894.260000 0.000000 1898.440000 0.630000 ;
      RECT 1889.660000 0.000000 1893.840000 0.630000 ;
      RECT 1885.520000 0.000000 1889.240000 0.630000 ;
      RECT 1880.920000 0.000000 1885.100000 0.630000 ;
      RECT 1876.320000 0.000000 1880.500000 0.630000 ;
      RECT 1871.720000 0.000000 1875.900000 0.630000 ;
      RECT 1867.120000 0.000000 1871.300000 0.630000 ;
      RECT 1862.520000 0.000000 1866.700000 0.630000 ;
      RECT 1857.920000 0.000000 1862.100000 0.630000 ;
      RECT 1853.320000 0.000000 1857.500000 0.630000 ;
      RECT 1849.180000 0.000000 1852.900000 0.630000 ;
      RECT 1844.580000 0.000000 1848.760000 0.630000 ;
      RECT 1839.980000 0.000000 1844.160000 0.630000 ;
      RECT 1835.380000 0.000000 1839.560000 0.630000 ;
      RECT 1830.780000 0.000000 1834.960000 0.630000 ;
      RECT 1826.180000 0.000000 1830.360000 0.630000 ;
      RECT 1821.580000 0.000000 1825.760000 0.630000 ;
      RECT 1816.980000 0.000000 1821.160000 0.630000 ;
      RECT 1812.840000 0.000000 1816.560000 0.630000 ;
      RECT 1808.240000 0.000000 1812.420000 0.630000 ;
      RECT 1803.640000 0.000000 1807.820000 0.630000 ;
      RECT 1799.040000 0.000000 1803.220000 0.630000 ;
      RECT 1794.440000 0.000000 1798.620000 0.630000 ;
      RECT 1789.840000 0.000000 1794.020000 0.630000 ;
      RECT 1785.240000 0.000000 1789.420000 0.630000 ;
      RECT 1780.640000 0.000000 1784.820000 0.630000 ;
      RECT 1776.500000 0.000000 1780.220000 0.630000 ;
      RECT 1771.900000 0.000000 1776.080000 0.630000 ;
      RECT 1767.300000 0.000000 1771.480000 0.630000 ;
      RECT 1762.700000 0.000000 1766.880000 0.630000 ;
      RECT 1758.100000 0.000000 1762.280000 0.630000 ;
      RECT 1753.500000 0.000000 1757.680000 0.630000 ;
      RECT 1748.900000 0.000000 1753.080000 0.630000 ;
      RECT 1744.300000 0.000000 1748.480000 0.630000 ;
      RECT 1740.160000 0.000000 1743.880000 0.630000 ;
      RECT 1735.560000 0.000000 1739.740000 0.630000 ;
      RECT 1730.960000 0.000000 1735.140000 0.630000 ;
      RECT 1726.360000 0.000000 1730.540000 0.630000 ;
      RECT 1721.760000 0.000000 1725.940000 0.630000 ;
      RECT 1717.160000 0.000000 1721.340000 0.630000 ;
      RECT 1712.560000 0.000000 1716.740000 0.630000 ;
      RECT 1707.960000 0.000000 1712.140000 0.630000 ;
      RECT 1703.820000 0.000000 1707.540000 0.630000 ;
      RECT 1699.220000 0.000000 1703.400000 0.630000 ;
      RECT 1694.620000 0.000000 1698.800000 0.630000 ;
      RECT 1690.020000 0.000000 1694.200000 0.630000 ;
      RECT 1685.420000 0.000000 1689.600000 0.630000 ;
      RECT 1680.820000 0.000000 1685.000000 0.630000 ;
      RECT 1676.220000 0.000000 1680.400000 0.630000 ;
      RECT 1671.620000 0.000000 1675.800000 0.630000 ;
      RECT 1667.480000 0.000000 1671.200000 0.630000 ;
      RECT 1662.880000 0.000000 1667.060000 0.630000 ;
      RECT 1658.280000 0.000000 1662.460000 0.630000 ;
      RECT 1653.680000 0.000000 1657.860000 0.630000 ;
      RECT 1649.080000 0.000000 1653.260000 0.630000 ;
      RECT 1644.480000 0.000000 1648.660000 0.630000 ;
      RECT 1639.880000 0.000000 1644.060000 0.630000 ;
      RECT 1635.280000 0.000000 1639.460000 0.630000 ;
      RECT 1631.140000 0.000000 1634.860000 0.630000 ;
      RECT 1626.540000 0.000000 1630.720000 0.630000 ;
      RECT 1621.940000 0.000000 1626.120000 0.630000 ;
      RECT 1617.340000 0.000000 1621.520000 0.630000 ;
      RECT 1612.740000 0.000000 1616.920000 0.630000 ;
      RECT 1608.140000 0.000000 1612.320000 0.630000 ;
      RECT 1603.540000 0.000000 1607.720000 0.630000 ;
      RECT 1598.940000 0.000000 1603.120000 0.630000 ;
      RECT 1594.800000 0.000000 1598.520000 0.630000 ;
      RECT 1590.200000 0.000000 1594.380000 0.630000 ;
      RECT 1585.600000 0.000000 1589.780000 0.630000 ;
      RECT 1581.000000 0.000000 1585.180000 0.630000 ;
      RECT 1576.400000 0.000000 1580.580000 0.630000 ;
      RECT 1571.800000 0.000000 1575.980000 0.630000 ;
      RECT 1567.200000 0.000000 1571.380000 0.630000 ;
      RECT 1562.600000 0.000000 1566.780000 0.630000 ;
      RECT 1558.460000 0.000000 1562.180000 0.630000 ;
      RECT 1553.860000 0.000000 1558.040000 0.630000 ;
      RECT 1549.260000 0.000000 1553.440000 0.630000 ;
      RECT 1544.660000 0.000000 1548.840000 0.630000 ;
      RECT 1540.060000 0.000000 1544.240000 0.630000 ;
      RECT 1535.460000 0.000000 1539.640000 0.630000 ;
      RECT 1530.860000 0.000000 1535.040000 0.630000 ;
      RECT 1526.260000 0.000000 1530.440000 0.630000 ;
      RECT 1521.660000 0.000000 1525.840000 0.630000 ;
      RECT 1517.520000 0.000000 1521.240000 0.630000 ;
      RECT 1512.920000 0.000000 1517.100000 0.630000 ;
      RECT 1508.320000 0.000000 1512.500000 0.630000 ;
      RECT 1503.720000 0.000000 1507.900000 0.630000 ;
      RECT 1499.120000 0.000000 1503.300000 0.630000 ;
      RECT 1494.520000 0.000000 1498.700000 0.630000 ;
      RECT 1489.920000 0.000000 1494.100000 0.630000 ;
      RECT 1485.320000 0.000000 1489.500000 0.630000 ;
      RECT 1481.180000 0.000000 1484.900000 0.630000 ;
      RECT 1476.580000 0.000000 1480.760000 0.630000 ;
      RECT 1471.980000 0.000000 1476.160000 0.630000 ;
      RECT 1467.380000 0.000000 1471.560000 0.630000 ;
      RECT 1462.780000 0.000000 1466.960000 0.630000 ;
      RECT 1458.180000 0.000000 1462.360000 0.630000 ;
      RECT 1453.580000 0.000000 1457.760000 0.630000 ;
      RECT 1448.980000 0.000000 1453.160000 0.630000 ;
      RECT 1444.840000 0.000000 1448.560000 0.630000 ;
      RECT 1440.240000 0.000000 1444.420000 0.630000 ;
      RECT 1435.640000 0.000000 1439.820000 0.630000 ;
      RECT 1431.040000 0.000000 1435.220000 0.630000 ;
      RECT 1426.440000 0.000000 1430.620000 0.630000 ;
      RECT 1421.840000 0.000000 1426.020000 0.630000 ;
      RECT 1417.240000 0.000000 1421.420000 0.630000 ;
      RECT 1412.640000 0.000000 1416.820000 0.630000 ;
      RECT 1408.500000 0.000000 1412.220000 0.630000 ;
      RECT 1403.900000 0.000000 1408.080000 0.630000 ;
      RECT 1399.300000 0.000000 1403.480000 0.630000 ;
      RECT 1394.700000 0.000000 1398.880000 0.630000 ;
      RECT 1390.100000 0.000000 1394.280000 0.630000 ;
      RECT 1385.500000 0.000000 1389.680000 0.630000 ;
      RECT 1380.900000 0.000000 1385.080000 0.630000 ;
      RECT 1376.300000 0.000000 1380.480000 0.630000 ;
      RECT 1372.160000 0.000000 1375.880000 0.630000 ;
      RECT 1367.560000 0.000000 1371.740000 0.630000 ;
      RECT 1362.960000 0.000000 1367.140000 0.630000 ;
      RECT 1358.360000 0.000000 1362.540000 0.630000 ;
      RECT 1353.760000 0.000000 1357.940000 0.630000 ;
      RECT 1349.160000 0.000000 1353.340000 0.630000 ;
      RECT 1344.560000 0.000000 1348.740000 0.630000 ;
      RECT 1339.960000 0.000000 1344.140000 0.630000 ;
      RECT 1335.820000 0.000000 1339.540000 0.630000 ;
      RECT 1331.220000 0.000000 1335.400000 0.630000 ;
      RECT 1326.620000 0.000000 1330.800000 0.630000 ;
      RECT 1322.020000 0.000000 1326.200000 0.630000 ;
      RECT 1317.420000 0.000000 1321.600000 0.630000 ;
      RECT 1312.820000 0.000000 1317.000000 0.630000 ;
      RECT 1308.220000 0.000000 1312.400000 0.630000 ;
      RECT 1303.620000 0.000000 1307.800000 0.630000 ;
      RECT 1299.480000 0.000000 1303.200000 0.630000 ;
      RECT 1294.880000 0.000000 1299.060000 0.630000 ;
      RECT 1290.280000 0.000000 1294.460000 0.630000 ;
      RECT 1285.680000 0.000000 1289.860000 0.630000 ;
      RECT 1281.080000 0.000000 1285.260000 0.630000 ;
      RECT 1276.480000 0.000000 1280.660000 0.630000 ;
      RECT 1271.880000 0.000000 1276.060000 0.630000 ;
      RECT 1267.280000 0.000000 1271.460000 0.630000 ;
      RECT 1263.140000 0.000000 1266.860000 0.630000 ;
      RECT 1258.540000 0.000000 1262.720000 0.630000 ;
      RECT 1253.940000 0.000000 1258.120000 0.630000 ;
      RECT 1249.340000 0.000000 1253.520000 0.630000 ;
      RECT 1244.740000 0.000000 1248.920000 0.630000 ;
      RECT 1240.140000 0.000000 1244.320000 0.630000 ;
      RECT 1235.540000 0.000000 1239.720000 0.630000 ;
      RECT 1230.940000 0.000000 1235.120000 0.630000 ;
      RECT 1226.800000 0.000000 1230.520000 0.630000 ;
      RECT 1222.200000 0.000000 1226.380000 0.630000 ;
      RECT 1217.600000 0.000000 1221.780000 0.630000 ;
      RECT 1213.000000 0.000000 1217.180000 0.630000 ;
      RECT 1208.400000 0.000000 1212.580000 0.630000 ;
      RECT 1203.800000 0.000000 1207.980000 0.630000 ;
      RECT 1199.200000 0.000000 1203.380000 0.630000 ;
      RECT 1194.600000 0.000000 1198.780000 0.630000 ;
      RECT 1190.460000 0.000000 1194.180000 0.630000 ;
      RECT 1185.860000 0.000000 1190.040000 0.630000 ;
      RECT 1181.260000 0.000000 1185.440000 0.630000 ;
      RECT 1176.660000 0.000000 1180.840000 0.630000 ;
      RECT 1172.060000 0.000000 1176.240000 0.630000 ;
      RECT 1167.460000 0.000000 1171.640000 0.630000 ;
      RECT 1162.860000 0.000000 1167.040000 0.630000 ;
      RECT 1158.260000 0.000000 1162.440000 0.630000 ;
      RECT 1154.120000 0.000000 1157.840000 0.630000 ;
      RECT 1149.520000 0.000000 1153.700000 0.630000 ;
      RECT 1144.920000 0.000000 1149.100000 0.630000 ;
      RECT 1140.320000 0.000000 1144.500000 0.630000 ;
      RECT 1135.720000 0.000000 1139.900000 0.630000 ;
      RECT 1131.120000 0.000000 1135.300000 0.630000 ;
      RECT 1126.520000 0.000000 1130.700000 0.630000 ;
      RECT 1121.920000 0.000000 1126.100000 0.630000 ;
      RECT 1117.780000 0.000000 1121.500000 0.630000 ;
      RECT 1113.180000 0.000000 1117.360000 0.630000 ;
      RECT 1108.580000 0.000000 1112.760000 0.630000 ;
      RECT 1103.980000 0.000000 1108.160000 0.630000 ;
      RECT 1099.380000 0.000000 1103.560000 0.630000 ;
      RECT 1094.780000 0.000000 1098.960000 0.630000 ;
      RECT 1090.180000 0.000000 1094.360000 0.630000 ;
      RECT 1085.580000 0.000000 1089.760000 0.630000 ;
      RECT 1081.440000 0.000000 1085.160000 0.630000 ;
      RECT 1076.840000 0.000000 1081.020000 0.630000 ;
      RECT 1072.240000 0.000000 1076.420000 0.630000 ;
      RECT 1067.640000 0.000000 1071.820000 0.630000 ;
      RECT 1063.040000 0.000000 1067.220000 0.630000 ;
      RECT 1058.440000 0.000000 1062.620000 0.630000 ;
      RECT 1053.840000 0.000000 1058.020000 0.630000 ;
      RECT 1049.240000 0.000000 1053.420000 0.630000 ;
      RECT 1045.100000 0.000000 1048.820000 0.630000 ;
      RECT 1040.500000 0.000000 1044.680000 0.630000 ;
      RECT 1035.900000 0.000000 1040.080000 0.630000 ;
      RECT 1031.300000 0.000000 1035.480000 0.630000 ;
      RECT 1026.700000 0.000000 1030.880000 0.630000 ;
      RECT 1022.100000 0.000000 1026.280000 0.630000 ;
      RECT 1017.500000 0.000000 1021.680000 0.630000 ;
      RECT 1012.900000 0.000000 1017.080000 0.630000 ;
      RECT 1008.300000 0.000000 1012.480000 0.630000 ;
      RECT 1004.160000 0.000000 1007.880000 0.630000 ;
      RECT 999.560000 0.000000 1003.740000 0.630000 ;
      RECT 994.960000 0.000000 999.140000 0.630000 ;
      RECT 990.360000 0.000000 994.540000 0.630000 ;
      RECT 985.760000 0.000000 989.940000 0.630000 ;
      RECT 981.160000 0.000000 985.340000 0.630000 ;
      RECT 976.560000 0.000000 980.740000 0.630000 ;
      RECT 971.960000 0.000000 976.140000 0.630000 ;
      RECT 967.820000 0.000000 971.540000 0.630000 ;
      RECT 963.220000 0.000000 967.400000 0.630000 ;
      RECT 958.620000 0.000000 962.800000 0.630000 ;
      RECT 954.020000 0.000000 958.200000 0.630000 ;
      RECT 949.420000 0.000000 953.600000 0.630000 ;
      RECT 944.820000 0.000000 949.000000 0.630000 ;
      RECT 940.220000 0.000000 944.400000 0.630000 ;
      RECT 935.620000 0.000000 939.800000 0.630000 ;
      RECT 931.480000 0.000000 935.200000 0.630000 ;
      RECT 926.880000 0.000000 931.060000 0.630000 ;
      RECT 922.280000 0.000000 926.460000 0.630000 ;
      RECT 917.680000 0.000000 921.860000 0.630000 ;
      RECT 913.080000 0.000000 917.260000 0.630000 ;
      RECT 908.480000 0.000000 912.660000 0.630000 ;
      RECT 903.880000 0.000000 908.060000 0.630000 ;
      RECT 899.280000 0.000000 903.460000 0.630000 ;
      RECT 895.140000 0.000000 898.860000 0.630000 ;
      RECT 890.540000 0.000000 894.720000 0.630000 ;
      RECT 885.940000 0.000000 890.120000 0.630000 ;
      RECT 881.340000 0.000000 885.520000 0.630000 ;
      RECT 876.740000 0.000000 880.920000 0.630000 ;
      RECT 872.140000 0.000000 876.320000 0.630000 ;
      RECT 867.540000 0.000000 871.720000 0.630000 ;
      RECT 862.940000 0.000000 867.120000 0.630000 ;
      RECT 858.800000 0.000000 862.520000 0.630000 ;
      RECT 854.200000 0.000000 858.380000 0.630000 ;
      RECT 849.600000 0.000000 853.780000 0.630000 ;
      RECT 845.000000 0.000000 849.180000 0.630000 ;
      RECT 840.400000 0.000000 844.580000 0.630000 ;
      RECT 835.800000 0.000000 839.980000 0.630000 ;
      RECT 831.200000 0.000000 835.380000 0.630000 ;
      RECT 826.600000 0.000000 830.780000 0.630000 ;
      RECT 822.460000 0.000000 826.180000 0.630000 ;
      RECT 817.860000 0.000000 822.040000 0.630000 ;
      RECT 813.260000 0.000000 817.440000 0.630000 ;
      RECT 808.660000 0.000000 812.840000 0.630000 ;
      RECT 804.060000 0.000000 808.240000 0.630000 ;
      RECT 799.460000 0.000000 803.640000 0.630000 ;
      RECT 794.860000 0.000000 799.040000 0.630000 ;
      RECT 790.260000 0.000000 794.440000 0.630000 ;
      RECT 786.120000 0.000000 789.840000 0.630000 ;
      RECT 781.520000 0.000000 785.700000 0.630000 ;
      RECT 776.920000 0.000000 781.100000 0.630000 ;
      RECT 772.320000 0.000000 776.500000 0.630000 ;
      RECT 767.720000 0.000000 771.900000 0.630000 ;
      RECT 763.120000 0.000000 767.300000 0.630000 ;
      RECT 758.520000 0.000000 762.700000 0.630000 ;
      RECT 753.920000 0.000000 758.100000 0.630000 ;
      RECT 749.780000 0.000000 753.500000 0.630000 ;
      RECT 745.180000 0.000000 749.360000 0.630000 ;
      RECT 740.580000 0.000000 744.760000 0.630000 ;
      RECT 735.980000 0.000000 740.160000 0.630000 ;
      RECT 731.380000 0.000000 735.560000 0.630000 ;
      RECT 726.780000 0.000000 730.960000 0.630000 ;
      RECT 722.180000 0.000000 726.360000 0.630000 ;
      RECT 717.580000 0.000000 721.760000 0.630000 ;
      RECT 713.440000 0.000000 717.160000 0.630000 ;
      RECT 708.840000 0.000000 713.020000 0.630000 ;
      RECT 704.240000 0.000000 708.420000 0.630000 ;
      RECT 699.640000 0.000000 703.820000 0.630000 ;
      RECT 695.040000 0.000000 699.220000 0.630000 ;
      RECT 690.440000 0.000000 694.620000 0.630000 ;
      RECT 685.840000 0.000000 690.020000 0.630000 ;
      RECT 681.240000 0.000000 685.420000 0.630000 ;
      RECT 677.100000 0.000000 680.820000 0.630000 ;
      RECT 672.500000 0.000000 676.680000 0.630000 ;
      RECT 667.900000 0.000000 672.080000 0.630000 ;
      RECT 663.300000 0.000000 667.480000 0.630000 ;
      RECT 658.700000 0.000000 662.880000 0.630000 ;
      RECT 654.100000 0.000000 658.280000 0.630000 ;
      RECT 649.500000 0.000000 653.680000 0.630000 ;
      RECT 644.900000 0.000000 649.080000 0.630000 ;
      RECT 640.760000 0.000000 644.480000 0.630000 ;
      RECT 636.160000 0.000000 640.340000 0.630000 ;
      RECT 631.560000 0.000000 635.740000 0.630000 ;
      RECT 626.960000 0.000000 631.140000 0.630000 ;
      RECT 622.360000 0.000000 626.540000 0.630000 ;
      RECT 617.760000 0.000000 621.940000 0.630000 ;
      RECT 613.160000 0.000000 617.340000 0.630000 ;
      RECT 608.560000 0.000000 612.740000 0.630000 ;
      RECT 604.420000 0.000000 608.140000 0.630000 ;
      RECT 599.820000 0.000000 604.000000 0.630000 ;
      RECT 595.220000 0.000000 599.400000 0.630000 ;
      RECT 590.620000 0.000000 594.800000 0.630000 ;
      RECT 586.020000 0.000000 590.200000 0.630000 ;
      RECT 581.420000 0.000000 585.600000 0.630000 ;
      RECT 576.820000 0.000000 581.000000 0.630000 ;
      RECT 572.220000 0.000000 576.400000 0.630000 ;
      RECT 568.080000 0.000000 571.800000 0.630000 ;
      RECT 563.480000 0.000000 567.660000 0.630000 ;
      RECT 558.880000 0.000000 563.060000 0.630000 ;
      RECT 554.280000 0.000000 558.460000 0.630000 ;
      RECT 549.680000 0.000000 553.860000 0.630000 ;
      RECT 545.080000 0.000000 549.260000 0.630000 ;
      RECT 540.480000 0.000000 544.660000 0.630000 ;
      RECT 535.880000 0.000000 540.060000 0.630000 ;
      RECT 531.740000 0.000000 535.460000 0.630000 ;
      RECT 527.140000 0.000000 531.320000 0.630000 ;
      RECT 522.540000 0.000000 526.720000 0.630000 ;
      RECT 517.940000 0.000000 522.120000 0.630000 ;
      RECT 513.340000 0.000000 517.520000 0.630000 ;
      RECT 508.740000 0.000000 512.920000 0.630000 ;
      RECT 504.140000 0.000000 508.320000 0.630000 ;
      RECT 499.540000 0.000000 503.720000 0.630000 ;
      RECT 494.940000 0.000000 499.120000 0.630000 ;
      RECT 490.800000 0.000000 494.520000 0.630000 ;
      RECT 486.200000 0.000000 490.380000 0.630000 ;
      RECT 481.600000 0.000000 485.780000 0.630000 ;
      RECT 5.040000 0.000000 481.180000 0.630000 ;
      RECT 4.580000 0.000000 4.620000 0.630000 ;
      RECT 0.000000 0.000000 4.160000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 2954.780000 2239.740000 2960.040000 ;
      RECT 0.000000 2953.880000 2238.640000 2954.780000 ;
      RECT 0.000000 2904.760000 2239.740000 2953.880000 ;
      RECT 1.100000 2903.860000 2239.740000 2904.760000 ;
      RECT 0.000000 2902.930000 2239.740000 2903.860000 ;
      RECT 0.000000 2902.030000 2238.640000 2902.930000 ;
      RECT 0.000000 2849.250000 2239.740000 2902.030000 ;
      RECT 1.100000 2848.350000 2239.740000 2849.250000 ;
      RECT 0.000000 2846.200000 2239.740000 2848.350000 ;
      RECT 0.000000 2845.300000 2238.640000 2846.200000 ;
      RECT 0.000000 2793.130000 2239.740000 2845.300000 ;
      RECT 1.100000 2792.230000 2239.740000 2793.130000 ;
      RECT 0.000000 2732.740000 2239.740000 2792.230000 ;
      RECT 0.000000 2731.840000 2238.640000 2732.740000 ;
      RECT 0.000000 2681.500000 2239.740000 2731.840000 ;
      RECT 1.100000 2680.600000 2239.740000 2681.500000 ;
      RECT 0.000000 2675.400000 2239.740000 2680.600000 ;
      RECT 0.000000 2674.500000 2238.640000 2675.400000 ;
      RECT 0.000000 2625.380000 2239.740000 2674.500000 ;
      RECT 1.100000 2624.480000 2239.740000 2625.380000 ;
      RECT 0.000000 2618.670000 2239.740000 2624.480000 ;
      RECT 0.000000 2617.770000 2238.640000 2618.670000 ;
      RECT 0.000000 2569.870000 2239.740000 2617.770000 ;
      RECT 1.100000 2568.970000 2239.740000 2569.870000 ;
      RECT 0.000000 2504.600000 2239.740000 2568.970000 ;
      RECT 0.000000 2503.700000 2238.640000 2504.600000 ;
      RECT 0.000000 2458.240000 2239.740000 2503.700000 ;
      RECT 1.100000 2457.340000 2239.740000 2458.240000 ;
      RECT 0.000000 2447.870000 2239.740000 2457.340000 ;
      RECT 0.000000 2446.970000 2238.640000 2447.870000 ;
      RECT 0.000000 2402.120000 2239.740000 2446.970000 ;
      RECT 1.100000 2401.220000 2239.740000 2402.120000 ;
      RECT 0.000000 2391.140000 2239.740000 2401.220000 ;
      RECT 0.000000 2390.240000 2238.640000 2391.140000 ;
      RECT 0.000000 2346.610000 2239.740000 2390.240000 ;
      RECT 1.100000 2345.710000 2239.740000 2346.610000 ;
      RECT 0.000000 2277.070000 2239.740000 2345.710000 ;
      RECT 0.000000 2276.170000 2238.640000 2277.070000 ;
      RECT 0.000000 2234.980000 2239.740000 2276.170000 ;
      RECT 1.100000 2234.080000 2239.740000 2234.980000 ;
      RECT 0.000000 2220.340000 2239.740000 2234.080000 ;
      RECT 0.000000 2219.440000 2238.640000 2220.340000 ;
      RECT 0.000000 2178.860000 2239.740000 2219.440000 ;
      RECT 1.100000 2177.960000 2239.740000 2178.860000 ;
      RECT 0.000000 2163.000000 2239.740000 2177.960000 ;
      RECT 0.000000 2162.100000 2238.640000 2163.000000 ;
      RECT 0.000000 2122.740000 2239.740000 2162.100000 ;
      RECT 1.100000 2121.840000 2239.740000 2122.740000 ;
      RECT 0.000000 2049.540000 2239.740000 2121.840000 ;
      RECT 0.000000 2048.640000 2238.640000 2049.540000 ;
      RECT 0.000000 2011.110000 2239.740000 2048.640000 ;
      RECT 1.100000 2010.210000 2239.740000 2011.110000 ;
      RECT 0.000000 1992.200000 2239.740000 2010.210000 ;
      RECT 0.000000 1991.300000 2238.640000 1992.200000 ;
      RECT 0.000000 1955.600000 2239.740000 1991.300000 ;
      RECT 1.100000 1954.700000 2239.740000 1955.600000 ;
      RECT 0.000000 1935.470000 2239.740000 1954.700000 ;
      RECT 0.000000 1934.570000 2238.640000 1935.470000 ;
      RECT 0.000000 1899.480000 2239.740000 1934.570000 ;
      RECT 1.100000 1898.580000 2239.740000 1899.480000 ;
      RECT 0.000000 1821.400000 2239.740000 1898.580000 ;
      RECT 0.000000 1820.500000 2238.640000 1821.400000 ;
      RECT 0.000000 1787.850000 2239.740000 1820.500000 ;
      RECT 1.100000 1786.950000 2239.740000 1787.850000 ;
      RECT 0.000000 1764.670000 2239.740000 1786.950000 ;
      RECT 0.000000 1763.770000 2238.640000 1764.670000 ;
      RECT 0.000000 1732.340000 2239.740000 1763.770000 ;
      RECT 1.100000 1731.440000 2239.740000 1732.340000 ;
      RECT 0.000000 1707.940000 2239.740000 1731.440000 ;
      RECT 0.000000 1707.040000 2238.640000 1707.940000 ;
      RECT 0.000000 1676.220000 2239.740000 1707.040000 ;
      RECT 1.100000 1675.320000 2239.740000 1676.220000 ;
      RECT 0.000000 1593.870000 2239.740000 1675.320000 ;
      RECT 0.000000 1592.970000 2238.640000 1593.870000 ;
      RECT 0.000000 1564.590000 2239.740000 1592.970000 ;
      RECT 1.100000 1563.690000 2239.740000 1564.590000 ;
      RECT 0.000000 1537.140000 2239.740000 1563.690000 ;
      RECT 0.000000 1536.240000 2238.640000 1537.140000 ;
      RECT 0.000000 1508.470000 2239.740000 1536.240000 ;
      RECT 1.100000 1507.570000 2239.740000 1508.470000 ;
      RECT 0.000000 1480.410000 2239.740000 1507.570000 ;
      RECT 0.000000 1479.510000 2238.640000 1480.410000 ;
      RECT 0.000000 1452.960000 2239.740000 1479.510000 ;
      RECT 1.100000 1452.060000 2239.740000 1452.960000 ;
      RECT 0.000000 1366.340000 2239.740000 1452.060000 ;
      RECT 0.000000 1365.440000 2238.640000 1366.340000 ;
      RECT 0.000000 1341.330000 2239.740000 1365.440000 ;
      RECT 1.100000 1340.430000 2239.740000 1341.330000 ;
      RECT 0.000000 1309.610000 2239.740000 1340.430000 ;
      RECT 0.000000 1308.710000 2238.640000 1309.610000 ;
      RECT 0.000000 1285.210000 2239.740000 1308.710000 ;
      RECT 1.100000 1284.310000 2239.740000 1285.210000 ;
      RECT 0.000000 1252.270000 2239.740000 1284.310000 ;
      RECT 0.000000 1251.370000 2238.640000 1252.270000 ;
      RECT 0.000000 1229.700000 2239.740000 1251.370000 ;
      RECT 1.100000 1228.800000 2239.740000 1229.700000 ;
      RECT 0.000000 1138.810000 2239.740000 1228.800000 ;
      RECT 0.000000 1137.910000 2238.640000 1138.810000 ;
      RECT 0.000000 1117.460000 2239.740000 1137.910000 ;
      RECT 1.100000 1116.560000 2239.740000 1117.460000 ;
      RECT 0.000000 1081.470000 2239.740000 1116.560000 ;
      RECT 0.000000 1080.570000 2238.640000 1081.470000 ;
      RECT 0.000000 1061.950000 2239.740000 1080.570000 ;
      RECT 1.100000 1061.050000 2239.740000 1061.950000 ;
      RECT 0.000000 1024.740000 2239.740000 1061.050000 ;
      RECT 0.000000 1023.840000 2238.640000 1024.740000 ;
      RECT 0.000000 1005.830000 2239.740000 1023.840000 ;
      RECT 1.100000 1004.930000 2239.740000 1005.830000 ;
      RECT 0.000000 968.010000 2239.740000 1004.930000 ;
      RECT 0.000000 967.110000 2238.640000 968.010000 ;
      RECT 0.000000 910.670000 2239.740000 967.110000 ;
      RECT 0.000000 909.770000 2238.640000 910.670000 ;
      RECT 0.000000 894.200000 2239.740000 909.770000 ;
      RECT 1.100000 893.300000 2239.740000 894.200000 ;
      RECT 0.000000 853.940000 2239.740000 893.300000 ;
      RECT 0.000000 853.040000 2238.640000 853.940000 ;
      RECT 0.000000 838.690000 2239.740000 853.040000 ;
      RECT 1.100000 837.790000 2239.740000 838.690000 ;
      RECT 0.000000 797.210000 2239.740000 837.790000 ;
      RECT 0.000000 796.310000 2238.640000 797.210000 ;
      RECT 0.000000 782.570000 2239.740000 796.310000 ;
      RECT 1.100000 781.670000 2239.740000 782.570000 ;
      RECT 0.000000 739.870000 2239.740000 781.670000 ;
      RECT 0.000000 738.970000 2238.640000 739.870000 ;
      RECT 0.000000 683.140000 2239.740000 738.970000 ;
      RECT 0.000000 682.240000 2238.640000 683.140000 ;
      RECT 0.000000 670.940000 2239.740000 682.240000 ;
      RECT 1.100000 670.040000 2239.740000 670.940000 ;
      RECT 0.000000 626.410000 2239.740000 670.040000 ;
      RECT 0.000000 625.510000 2238.640000 626.410000 ;
      RECT 0.000000 614.820000 2239.740000 625.510000 ;
      RECT 1.100000 613.920000 2239.740000 614.820000 ;
      RECT 0.000000 569.680000 2239.740000 613.920000 ;
      RECT 0.000000 568.780000 2238.640000 569.680000 ;
      RECT 0.000000 559.310000 2239.740000 568.780000 ;
      RECT 1.100000 558.410000 2239.740000 559.310000 ;
      RECT 0.000000 512.340000 2239.740000 558.410000 ;
      RECT 0.000000 511.440000 2238.640000 512.340000 ;
      RECT 0.000000 455.610000 2239.740000 511.440000 ;
      RECT 0.000000 454.710000 2238.640000 455.610000 ;
      RECT 0.000000 447.680000 2239.740000 454.710000 ;
      RECT 1.100000 446.780000 2239.740000 447.680000 ;
      RECT 0.000000 398.880000 2239.740000 446.780000 ;
      RECT 0.000000 397.980000 2238.640000 398.880000 ;
      RECT 0.000000 391.560000 2239.740000 397.980000 ;
      RECT 1.100000 390.660000 2239.740000 391.560000 ;
      RECT 0.000000 341.540000 2239.740000 390.660000 ;
      RECT 0.000000 340.640000 2238.640000 341.540000 ;
      RECT 0.000000 336.050000 2239.740000 340.640000 ;
      RECT 1.100000 335.150000 2239.740000 336.050000 ;
      RECT 0.000000 284.810000 2239.740000 335.150000 ;
      RECT 0.000000 283.910000 2238.640000 284.810000 ;
      RECT 0.000000 279.930000 2239.740000 283.910000 ;
      RECT 1.100000 279.030000 2239.740000 279.930000 ;
      RECT 0.000000 228.080000 2239.740000 279.030000 ;
      RECT 0.000000 227.180000 2238.640000 228.080000 ;
      RECT 0.000000 224.420000 2239.740000 227.180000 ;
      RECT 1.100000 223.520000 2239.740000 224.420000 ;
      RECT 0.000000 170.740000 2239.740000 223.520000 ;
      RECT 0.000000 169.840000 2238.640000 170.740000 ;
      RECT 0.000000 168.300000 2239.740000 169.840000 ;
      RECT 1.100000 167.400000 2239.740000 168.300000 ;
      RECT 0.000000 114.010000 2239.740000 167.400000 ;
      RECT 0.000000 113.110000 2238.640000 114.010000 ;
      RECT 0.000000 112.180000 2239.740000 113.110000 ;
      RECT 1.100000 111.280000 2239.740000 112.180000 ;
      RECT 0.000000 57.280000 2239.740000 111.280000 ;
      RECT 0.000000 56.670000 2238.640000 57.280000 ;
      RECT 1.100000 56.380000 2238.640000 56.670000 ;
      RECT 1.100000 55.770000 2239.740000 56.380000 ;
      RECT 0.000000 6.040000 2239.740000 55.770000 ;
      RECT 1.100000 5.140000 2239.740000 6.040000 ;
      RECT 0.000000 4.820000 2239.740000 5.140000 ;
      RECT 0.000000 3.920000 2238.640000 4.820000 ;
      RECT 0.000000 0.000000 2239.740000 3.920000 ;
    LAYER met4 ;
      RECT 0.000000 2955.630000 2239.740000 2960.040000 ;
      RECT 9.390000 2948.830000 2230.350000 2955.630000 ;
      RECT 2229.350000 10.530000 2230.350000 2948.830000 ;
      RECT 16.190000 10.530000 2223.550000 2948.830000 ;
      RECT 9.390000 10.530000 10.390000 2948.830000 ;
      RECT 2236.150000 3.730000 2239.740000 2955.630000 ;
      RECT 9.390000 3.730000 2230.350000 10.530000 ;
      RECT 0.000000 3.730000 3.590000 2955.630000 ;
      RECT 0.000000 0.000000 2239.740000 3.730000 ;
  END
END Ibtida_top_dffram_cv

END LIBRARY
