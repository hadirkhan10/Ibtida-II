##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sat Nov 27 17:36:59 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Ibtida_top_dffram_cv
  CLASS BLOCK ;
  SIZE 1742.480000 BY 1753.040000 ;
  FOREIGN Ibtida_top_dffram_cv 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300000 0.000000 4.440000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.160000 0.000000 0.300000 0.490000 ;
    END
  END wb_rst_i
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.440000 0.000000 583.580000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.300000 0.000000 579.440000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.700000 0.000000 574.840000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.100000 0.000000 570.240000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.500000 0.000000 565.640000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.900000 0.000000 561.040000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.300000 0.000000 556.440000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.160000 0.000000 552.300000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.560000 0.000000 547.700000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.960000 0.000000 543.100000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.360000 0.000000 538.500000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.760000 0.000000 533.900000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.160000 0.000000 529.300000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.020000 0.000000 525.160000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.420000 0.000000 520.560000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.820000 0.000000 515.960000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.220000 0.000000 511.360000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.620000 0.000000 506.760000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.020000 0.000000 502.160000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.880000 0.000000 498.020000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.280000 0.000000 493.420000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.680000 0.000000 488.820000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.080000 0.000000 484.220000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.480000 0.000000 479.620000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.880000 0.000000 475.020000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.280000 0.000000 470.420000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.140000 0.000000 466.280000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.540000 0.000000 461.680000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.940000 0.000000 457.080000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.340000 0.000000 452.480000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.740000 0.000000 447.880000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.140000 0.000000 443.280000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.000000 0.000000 439.140000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.400000 0.000000 434.540000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.800000 0.000000 429.940000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.200000 0.000000 425.340000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.600000 0.000000 420.740000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.000000 0.000000 416.140000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.860000 0.000000 412.000000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.260000 0.000000 407.400000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.660000 0.000000 402.800000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.060000 0.000000 398.200000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.460000 0.000000 393.600000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.860000 0.000000 389.000000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.720000 0.000000 384.860000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.120000 0.000000 380.260000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.520000 0.000000 375.660000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.920000 0.000000 371.060000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.320000 0.000000 366.460000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.720000 0.000000 361.860000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.580000 0.000000 357.720000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.980000 0.000000 353.120000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.380000 0.000000 348.520000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.780000 0.000000 343.920000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.180000 0.000000 339.320000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.580000 0.000000 334.720000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.440000 0.000000 330.580000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.840000 0.000000 325.980000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.240000 0.000000 321.380000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.640000 0.000000 316.780000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.040000 0.000000 312.180000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.440000 0.000000 307.580000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.300000 0.000000 303.440000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.700000 0.000000 298.840000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.100000 0.000000 294.240000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.500000 0.000000 289.640000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.900000 0.000000 285.040000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.300000 0.000000 280.440000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.160000 0.000000 276.300000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.560000 0.000000 271.700000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.960000 0.000000 267.100000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.360000 0.000000 262.500000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.760000 0.000000 257.900000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.160000 0.000000 253.300000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.560000 0.000000 248.700000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.420000 0.000000 244.560000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.820000 0.000000 239.960000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.220000 0.000000 235.360000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.620000 0.000000 230.760000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.020000 0.000000 226.160000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.420000 0.000000 221.560000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280000 0.000000 217.420000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680000 0.000000 212.820000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.080000 0.000000 208.220000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480000 0.000000 203.620000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.880000 0.000000 199.020000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.280000 0.000000 194.420000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.140000 0.000000 190.280000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.540000 0.000000 185.680000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940000 0.000000 181.080000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.340000 0.000000 176.480000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.740000 0.000000 171.880000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.140000 0.000000 167.280000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.000000 0.000000 163.140000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400000 0.000000 158.540000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.800000 0.000000 153.940000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.200000 0.000000 149.340000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.600000 0.000000 144.740000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.000000 0.000000 140.140000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.860000 0.000000 136.000000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.260000 0.000000 131.400000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.660000 0.000000 126.800000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.060000 0.000000 122.200000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460000 0.000000 117.600000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860000 0.000000 113.000000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.720000 0.000000 108.860000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120000 0.000000 104.260000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520000 0.000000 99.660000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920000 0.000000 95.060000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320000 0.000000 90.460000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.720000 0.000000 85.860000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.580000 0.000000 81.720000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980000 0.000000 77.120000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380000 0.000000 72.520000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.780000 0.000000 67.920000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180000 0.000000 63.320000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.580000 0.000000 58.720000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.440000 0.000000 54.580000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.840000 0.000000 49.980000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240000 0.000000 45.380000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640000 0.000000 40.780000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040000 0.000000 36.180000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.440000 0.000000 31.580000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300000 0.000000 27.440000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.700000 0.000000 22.840000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100000 0.000000 18.240000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.500000 0.000000 13.640000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900000 0.000000 9.040000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.580000 0.000000 1162.720000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.440000 0.000000 1158.580000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.840000 0.000000 1153.980000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.240000 0.000000 1149.380000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.640000 0.000000 1144.780000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.040000 0.000000 1140.180000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.440000 0.000000 1135.580000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.300000 0.000000 1131.440000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.700000 0.000000 1126.840000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.100000 0.000000 1122.240000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.500000 0.000000 1117.640000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.900000 0.000000 1113.040000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.300000 0.000000 1108.440000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.160000 0.000000 1104.300000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.560000 0.000000 1099.700000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.960000 0.000000 1095.100000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.360000 0.000000 1090.500000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.760000 0.000000 1085.900000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.160000 0.000000 1081.300000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.020000 0.000000 1077.160000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.420000 0.000000 1072.560000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.820000 0.000000 1067.960000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.220000 0.000000 1063.360000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.620000 0.000000 1058.760000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.020000 0.000000 1054.160000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.880000 0.000000 1050.020000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.280000 0.000000 1045.420000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.680000 0.000000 1040.820000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.080000 0.000000 1036.220000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.480000 0.000000 1031.620000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.880000 0.000000 1027.020000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.740000 0.000000 1022.880000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.140000 0.000000 1018.280000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.540000 0.000000 1013.680000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.940000 0.000000 1009.080000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.340000 0.000000 1004.480000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.740000 0.000000 999.880000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.140000 0.000000 995.280000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.000000 0.000000 991.140000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.400000 0.000000 986.540000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.800000 0.000000 981.940000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.200000 0.000000 977.340000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.600000 0.000000 972.740000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.000000 0.000000 968.140000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.860000 0.000000 964.000000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.260000 0.000000 959.400000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.660000 0.000000 954.800000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.060000 0.000000 950.200000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.460000 0.000000 945.600000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.860000 0.000000 941.000000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.720000 0.000000 936.860000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.120000 0.000000 932.260000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.520000 0.000000 927.660000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.920000 0.000000 923.060000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.320000 0.000000 918.460000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.720000 0.000000 913.860000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.580000 0.000000 909.720000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.980000 0.000000 905.120000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.380000 0.000000 900.520000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.780000 0.000000 895.920000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.180000 0.000000 891.320000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.580000 0.000000 886.720000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.440000 0.000000 882.580000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.840000 0.000000 877.980000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.240000 0.000000 873.380000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.640000 0.000000 868.780000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.040000 0.000000 864.180000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.440000 0.000000 859.580000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.300000 0.000000 855.440000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.700000 0.000000 850.840000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.100000 0.000000 846.240000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.500000 0.000000 841.640000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.900000 0.000000 837.040000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.300000 0.000000 832.440000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.160000 0.000000 828.300000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.560000 0.000000 823.700000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.960000 0.000000 819.100000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.360000 0.000000 814.500000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.760000 0.000000 809.900000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.160000 0.000000 805.300000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.020000 0.000000 801.160000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.420000 0.000000 796.560000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.820000 0.000000 791.960000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.220000 0.000000 787.360000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.620000 0.000000 782.760000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.020000 0.000000 778.160000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.880000 0.000000 774.020000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.280000 0.000000 769.420000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.680000 0.000000 764.820000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.080000 0.000000 760.220000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.480000 0.000000 755.620000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.880000 0.000000 751.020000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.280000 0.000000 746.420000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.140000 0.000000 742.280000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.540000 0.000000 737.680000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.940000 0.000000 733.080000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.340000 0.000000 728.480000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.740000 0.000000 723.880000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.140000 0.000000 719.280000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.000000 0.000000 715.140000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.400000 0.000000 710.540000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.800000 0.000000 705.940000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.200000 0.000000 701.340000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.600000 0.000000 696.740000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.000000 0.000000 692.140000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.860000 0.000000 688.000000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.260000 0.000000 683.400000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.660000 0.000000 678.800000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.060000 0.000000 674.200000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.460000 0.000000 669.600000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.860000 0.000000 665.000000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.720000 0.000000 660.860000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.120000 0.000000 656.260000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.520000 0.000000 651.660000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.920000 0.000000 647.060000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.320000 0.000000 642.460000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.720000 0.000000 637.860000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.580000 0.000000 633.720000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.980000 0.000000 629.120000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.380000 0.000000 624.520000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.780000 0.000000 619.920000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.180000 0.000000 615.320000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.580000 0.000000 610.720000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.440000 0.000000 606.580000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.840000 0.000000 601.980000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.240000 0.000000 597.380000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.640000 0.000000 592.780000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.040000 0.000000 588.180000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.180000 0.000000 1742.320000 0.490000 ;
    END
  END la_oen[127]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.580000 0.000000 1737.720000 0.490000 ;
    END
  END la_oen[126]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.980000 0.000000 1733.120000 0.490000 ;
    END
  END la_oen[125]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.380000 0.000000 1728.520000 0.490000 ;
    END
  END la_oen[124]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.780000 0.000000 1723.920000 0.490000 ;
    END
  END la_oen[123]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.180000 0.000000 1719.320000 0.490000 ;
    END
  END la_oen[122]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.580000 0.000000 1714.720000 0.490000 ;
    END
  END la_oen[121]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.440000 0.000000 1710.580000 0.490000 ;
    END
  END la_oen[120]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.840000 0.000000 1705.980000 0.490000 ;
    END
  END la_oen[119]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.240000 0.000000 1701.380000 0.490000 ;
    END
  END la_oen[118]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.640000 0.000000 1696.780000 0.490000 ;
    END
  END la_oen[117]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.040000 0.000000 1692.180000 0.490000 ;
    END
  END la_oen[116]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.440000 0.000000 1687.580000 0.490000 ;
    END
  END la_oen[115]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.300000 0.000000 1683.440000 0.490000 ;
    END
  END la_oen[114]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.700000 0.000000 1678.840000 0.490000 ;
    END
  END la_oen[113]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.100000 0.000000 1674.240000 0.490000 ;
    END
  END la_oen[112]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.500000 0.000000 1669.640000 0.490000 ;
    END
  END la_oen[111]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.900000 0.000000 1665.040000 0.490000 ;
    END
  END la_oen[110]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.300000 0.000000 1660.440000 0.490000 ;
    END
  END la_oen[109]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.160000 0.000000 1656.300000 0.490000 ;
    END
  END la_oen[108]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.560000 0.000000 1651.700000 0.490000 ;
    END
  END la_oen[107]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.960000 0.000000 1647.100000 0.490000 ;
    END
  END la_oen[106]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.360000 0.000000 1642.500000 0.490000 ;
    END
  END la_oen[105]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.760000 0.000000 1637.900000 0.490000 ;
    END
  END la_oen[104]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.160000 0.000000 1633.300000 0.490000 ;
    END
  END la_oen[103]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.020000 0.000000 1629.160000 0.490000 ;
    END
  END la_oen[102]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.420000 0.000000 1624.560000 0.490000 ;
    END
  END la_oen[101]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.820000 0.000000 1619.960000 0.490000 ;
    END
  END la_oen[100]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.220000 0.000000 1615.360000 0.490000 ;
    END
  END la_oen[99]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.620000 0.000000 1610.760000 0.490000 ;
    END
  END la_oen[98]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.020000 0.000000 1606.160000 0.490000 ;
    END
  END la_oen[97]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.880000 0.000000 1602.020000 0.490000 ;
    END
  END la_oen[96]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.280000 0.000000 1597.420000 0.490000 ;
    END
  END la_oen[95]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.680000 0.000000 1592.820000 0.490000 ;
    END
  END la_oen[94]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.080000 0.000000 1588.220000 0.490000 ;
    END
  END la_oen[93]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.480000 0.000000 1583.620000 0.490000 ;
    END
  END la_oen[92]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.880000 0.000000 1579.020000 0.490000 ;
    END
  END la_oen[91]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.740000 0.000000 1574.880000 0.490000 ;
    END
  END la_oen[90]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.140000 0.000000 1570.280000 0.490000 ;
    END
  END la_oen[89]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.540000 0.000000 1565.680000 0.490000 ;
    END
  END la_oen[88]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.940000 0.000000 1561.080000 0.490000 ;
    END
  END la_oen[87]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.340000 0.000000 1556.480000 0.490000 ;
    END
  END la_oen[86]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.740000 0.000000 1551.880000 0.490000 ;
    END
  END la_oen[85]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.600000 0.000000 1547.740000 0.490000 ;
    END
  END la_oen[84]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.000000 0.000000 1543.140000 0.490000 ;
    END
  END la_oen[83]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.400000 0.000000 1538.540000 0.490000 ;
    END
  END la_oen[82]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.800000 0.000000 1533.940000 0.490000 ;
    END
  END la_oen[81]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.200000 0.000000 1529.340000 0.490000 ;
    END
  END la_oen[80]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.600000 0.000000 1524.740000 0.490000 ;
    END
  END la_oen[79]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.460000 0.000000 1520.600000 0.490000 ;
    END
  END la_oen[78]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.860000 0.000000 1516.000000 0.490000 ;
    END
  END la_oen[77]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.260000 0.000000 1511.400000 0.490000 ;
    END
  END la_oen[76]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.660000 0.000000 1506.800000 0.490000 ;
    END
  END la_oen[75]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.060000 0.000000 1502.200000 0.490000 ;
    END
  END la_oen[74]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.460000 0.000000 1497.600000 0.490000 ;
    END
  END la_oen[73]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.320000 0.000000 1493.460000 0.490000 ;
    END
  END la_oen[72]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.720000 0.000000 1488.860000 0.490000 ;
    END
  END la_oen[71]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.120000 0.000000 1484.260000 0.490000 ;
    END
  END la_oen[70]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.520000 0.000000 1479.660000 0.490000 ;
    END
  END la_oen[69]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.920000 0.000000 1475.060000 0.490000 ;
    END
  END la_oen[68]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.320000 0.000000 1470.460000 0.490000 ;
    END
  END la_oen[67]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.720000 0.000000 1465.860000 0.490000 ;
    END
  END la_oen[66]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.580000 0.000000 1461.720000 0.490000 ;
    END
  END la_oen[65]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.980000 0.000000 1457.120000 0.490000 ;
    END
  END la_oen[64]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.380000 0.000000 1452.520000 0.490000 ;
    END
  END la_oen[63]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.780000 0.000000 1447.920000 0.490000 ;
    END
  END la_oen[62]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.180000 0.000000 1443.320000 0.490000 ;
    END
  END la_oen[61]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.580000 0.000000 1438.720000 0.490000 ;
    END
  END la_oen[60]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.440000 0.000000 1434.580000 0.490000 ;
    END
  END la_oen[59]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.840000 0.000000 1429.980000 0.490000 ;
    END
  END la_oen[58]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.240000 0.000000 1425.380000 0.490000 ;
    END
  END la_oen[57]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.640000 0.000000 1420.780000 0.490000 ;
    END
  END la_oen[56]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.040000 0.000000 1416.180000 0.490000 ;
    END
  END la_oen[55]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.440000 0.000000 1411.580000 0.490000 ;
    END
  END la_oen[54]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.300000 0.000000 1407.440000 0.490000 ;
    END
  END la_oen[53]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.700000 0.000000 1402.840000 0.490000 ;
    END
  END la_oen[52]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.100000 0.000000 1398.240000 0.490000 ;
    END
  END la_oen[51]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.500000 0.000000 1393.640000 0.490000 ;
    END
  END la_oen[50]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.900000 0.000000 1389.040000 0.490000 ;
    END
  END la_oen[49]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.300000 0.000000 1384.440000 0.490000 ;
    END
  END la_oen[48]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.160000 0.000000 1380.300000 0.490000 ;
    END
  END la_oen[47]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.560000 0.000000 1375.700000 0.490000 ;
    END
  END la_oen[46]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.960000 0.000000 1371.100000 0.490000 ;
    END
  END la_oen[45]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.360000 0.000000 1366.500000 0.490000 ;
    END
  END la_oen[44]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.760000 0.000000 1361.900000 0.490000 ;
    END
  END la_oen[43]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.160000 0.000000 1357.300000 0.490000 ;
    END
  END la_oen[42]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.020000 0.000000 1353.160000 0.490000 ;
    END
  END la_oen[41]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.420000 0.000000 1348.560000 0.490000 ;
    END
  END la_oen[40]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.820000 0.000000 1343.960000 0.490000 ;
    END
  END la_oen[39]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.220000 0.000000 1339.360000 0.490000 ;
    END
  END la_oen[38]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.620000 0.000000 1334.760000 0.490000 ;
    END
  END la_oen[37]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.020000 0.000000 1330.160000 0.490000 ;
    END
  END la_oen[36]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.880000 0.000000 1326.020000 0.490000 ;
    END
  END la_oen[35]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.280000 0.000000 1321.420000 0.490000 ;
    END
  END la_oen[34]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.680000 0.000000 1316.820000 0.490000 ;
    END
  END la_oen[33]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.080000 0.000000 1312.220000 0.490000 ;
    END
  END la_oen[32]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.480000 0.000000 1307.620000 0.490000 ;
    END
  END la_oen[31]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.880000 0.000000 1303.020000 0.490000 ;
    END
  END la_oen[30]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.740000 0.000000 1298.880000 0.490000 ;
    END
  END la_oen[29]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.140000 0.000000 1294.280000 0.490000 ;
    END
  END la_oen[28]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.540000 0.000000 1289.680000 0.490000 ;
    END
  END la_oen[27]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.940000 0.000000 1285.080000 0.490000 ;
    END
  END la_oen[26]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.340000 0.000000 1280.480000 0.490000 ;
    END
  END la_oen[25]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.740000 0.000000 1275.880000 0.490000 ;
    END
  END la_oen[24]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.600000 0.000000 1271.740000 0.490000 ;
    END
  END la_oen[23]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.000000 0.000000 1267.140000 0.490000 ;
    END
  END la_oen[22]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.400000 0.000000 1262.540000 0.490000 ;
    END
  END la_oen[21]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.800000 0.000000 1257.940000 0.490000 ;
    END
  END la_oen[20]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.200000 0.000000 1253.340000 0.490000 ;
    END
  END la_oen[19]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.600000 0.000000 1248.740000 0.490000 ;
    END
  END la_oen[18]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.460000 0.000000 1244.600000 0.490000 ;
    END
  END la_oen[17]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.860000 0.000000 1240.000000 0.490000 ;
    END
  END la_oen[16]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.260000 0.000000 1235.400000 0.490000 ;
    END
  END la_oen[15]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.660000 0.000000 1230.800000 0.490000 ;
    END
  END la_oen[14]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.060000 0.000000 1226.200000 0.490000 ;
    END
  END la_oen[13]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.460000 0.000000 1221.600000 0.490000 ;
    END
  END la_oen[12]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.860000 0.000000 1217.000000 0.490000 ;
    END
  END la_oen[11]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.720000 0.000000 1212.860000 0.490000 ;
    END
  END la_oen[10]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.120000 0.000000 1208.260000 0.490000 ;
    END
  END la_oen[9]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.520000 0.000000 1203.660000 0.490000 ;
    END
  END la_oen[8]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.920000 0.000000 1199.060000 0.490000 ;
    END
  END la_oen[7]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.320000 0.000000 1194.460000 0.490000 ;
    END
  END la_oen[6]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.720000 0.000000 1189.860000 0.490000 ;
    END
  END la_oen[5]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.580000 0.000000 1185.720000 0.490000 ;
    END
  END la_oen[4]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.980000 0.000000 1181.120000 0.490000 ;
    END
  END la_oen[3]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.380000 0.000000 1176.520000 0.490000 ;
    END
  END la_oen[2]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.780000 0.000000 1171.920000 0.490000 ;
    END
  END la_oen[1]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.180000 0.000000 1167.320000 0.490000 ;
    END
  END la_oen[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 85.960000 0.800000 86.260000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 214.060000 0.800000 214.360000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 342.160000 0.800000 342.460000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 470.260000 0.800000 470.560000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 598.360000 0.800000 598.660000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 726.460000 0.800000 726.760000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 854.560000 0.800000 854.860000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 983.270000 0.800000 983.570000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1111.370000 0.800000 1111.670000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1239.470000 0.800000 1239.770000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1367.570000 0.800000 1367.870000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1495.670000 0.800000 1495.970000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1623.770000 0.800000 1624.070000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1751.870000 0.800000 1752.170000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.020000 1752.550000 134.160000 1753.040000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.040000 1752.550000 335.180000 1753.040000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.060000 1752.550000 536.200000 1753.040000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.080000 1752.550000 737.220000 1753.040000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.100000 1752.550000 938.240000 1753.040000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.120000 1752.550000 1139.260000 1753.040000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.140000 1752.550000 1340.280000 1753.040000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.160000 1752.550000 1541.300000 1753.040000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.180000 1752.550000 1742.320000 1753.040000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1672.570000 1742.480000 1672.870000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1553.010000 1742.480000 1553.310000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1433.450000 1742.480000 1433.750000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1314.500000 1742.480000 1314.800000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1194.940000 1742.480000 1195.240000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1075.380000 1742.480000 1075.680000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 955.820000 1742.480000 956.120000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 836.260000 1742.480000 836.560000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 716.700000 1742.480000 717.000000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 597.750000 1742.480000 598.050000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 478.190000 1742.480000 478.490000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 358.630000 1742.480000 358.930000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 239.070000 1742.480000 239.370000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 119.510000 1742.480000 119.810000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 0.560000 1742.480000 0.860000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.260000 0.800000 43.560000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 171.360000 0.800000 171.660000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 299.460000 0.800000 299.760000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 427.560000 0.800000 427.860000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 555.660000 0.800000 555.960000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 683.760000 0.800000 684.060000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 811.860000 0.800000 812.160000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 940.570000 0.800000 940.870000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1068.670000 0.800000 1068.970000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1196.770000 0.800000 1197.070000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1324.870000 0.800000 1325.170000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1452.970000 0.800000 1453.270000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1581.070000 0.800000 1581.370000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1709.170000 0.800000 1709.470000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860000 1752.550000 67.000000 1753.040000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.880000 1752.550000 268.020000 1753.040000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.900000 1752.550000 469.040000 1753.040000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.920000 1752.550000 670.060000 1753.040000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.940000 1752.550000 871.080000 1753.040000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.960000 1752.550000 1072.100000 1753.040000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.980000 1752.550000 1273.120000 1753.040000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.000000 1752.550000 1474.140000 1753.040000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.020000 1752.550000 1675.160000 1753.040000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1712.220000 1742.480000 1712.520000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1592.660000 1742.480000 1592.960000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1473.710000 1742.480000 1474.010000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1354.150000 1742.480000 1354.450000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1234.590000 1742.480000 1234.890000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1115.030000 1742.480000 1115.330000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 995.470000 1742.480000 995.770000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 875.910000 1742.480000 876.210000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 756.960000 1742.480000 757.260000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 637.400000 1742.480000 637.700000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 517.840000 1742.480000 518.140000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 398.280000 1742.480000 398.580000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 278.720000 1742.480000 279.020000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 159.770000 1742.480000 160.070000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 40.210000 1742.480000 40.510000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.560000 0.800000 0.860000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.660000 0.800000 128.960000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 256.760000 0.800000 257.060000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 384.860000 0.800000 385.160000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 512.960000 0.800000 513.260000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 641.060000 0.800000 641.360000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 769.160000 0.800000 769.460000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 897.870000 0.800000 898.170000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1025.970000 0.800000 1026.270000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1154.070000 0.800000 1154.370000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1282.170000 0.800000 1282.470000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1410.270000 0.800000 1410.570000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1538.370000 0.800000 1538.670000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1666.470000 0.800000 1666.770000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.160000 1752.550000 0.300000 1753.040000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.720000 1752.550000 200.860000 1753.040000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.740000 1752.550000 401.880000 1753.040000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.760000 1752.550000 602.900000 1753.040000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.780000 1752.550000 803.920000 1753.040000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.800000 1752.550000 1004.940000 1753.040000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.820000 1752.550000 1205.960000 1753.040000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.840000 1752.550000 1406.980000 1753.040000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.860000 1752.550000 1608.000000 1753.040000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1752.480000 1742.480000 1752.780000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1632.920000 1742.480000 1633.220000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1513.360000 1742.480000 1513.660000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1393.800000 1742.480000 1394.100000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1274.240000 1742.480000 1274.540000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1154.680000 1742.480000 1154.980000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 1035.730000 1742.480000 1036.030000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 916.170000 1742.480000 916.470000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 796.610000 1742.480000 796.910000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 677.050000 1742.480000 677.350000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 557.490000 1742.480000 557.790000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 437.930000 1742.480000 438.230000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 318.980000 1742.480000 319.280000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 199.420000 1742.480000 199.720000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1741.680000 79.860000 1742.480000 80.160000 ;
    END
  END io_oeb[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1726.690000 10.930000 1731.690000 1741.090000 ;
    END
    PORT
      LAYER met4 ;
        RECT 10.790000 10.930000 15.790000 1741.090000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.990000 4.130000 8.990000 1747.890000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.490000 4.130000 1738.490000 1747.890000 ;
    END
  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1742.480000 1753.040000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1742.480000 1753.040000 ;
    LAYER met2 ;
      RECT 1742.460000 1752.410000 1742.480000 1753.040000 ;
      RECT 1675.300000 1752.410000 1742.040000 1753.040000 ;
      RECT 1608.140000 1752.410000 1674.880000 1753.040000 ;
      RECT 1541.440000 1752.410000 1607.720000 1753.040000 ;
      RECT 1474.280000 1752.410000 1541.020000 1753.040000 ;
      RECT 1407.120000 1752.410000 1473.860000 1753.040000 ;
      RECT 1340.420000 1752.410000 1406.700000 1753.040000 ;
      RECT 1273.260000 1752.410000 1340.000000 1753.040000 ;
      RECT 1206.100000 1752.410000 1272.840000 1753.040000 ;
      RECT 1139.400000 1752.410000 1205.680000 1753.040000 ;
      RECT 1072.240000 1752.410000 1138.980000 1753.040000 ;
      RECT 1005.080000 1752.410000 1071.820000 1753.040000 ;
      RECT 938.380000 1752.410000 1004.660000 1753.040000 ;
      RECT 871.220000 1752.410000 937.960000 1753.040000 ;
      RECT 804.060000 1752.410000 870.800000 1753.040000 ;
      RECT 737.360000 1752.410000 803.640000 1753.040000 ;
      RECT 670.200000 1752.410000 736.940000 1753.040000 ;
      RECT 603.040000 1752.410000 669.780000 1753.040000 ;
      RECT 536.340000 1752.410000 602.620000 1753.040000 ;
      RECT 469.180000 1752.410000 535.920000 1753.040000 ;
      RECT 402.020000 1752.410000 468.760000 1753.040000 ;
      RECT 335.320000 1752.410000 401.600000 1753.040000 ;
      RECT 268.160000 1752.410000 334.900000 1753.040000 ;
      RECT 201.000000 1752.410000 267.740000 1753.040000 ;
      RECT 134.300000 1752.410000 200.580000 1753.040000 ;
      RECT 67.140000 1752.410000 133.880000 1753.040000 ;
      RECT 0.440000 1752.410000 66.720000 1753.040000 ;
      RECT 0.000000 1752.410000 0.020000 1753.040000 ;
      RECT 0.000000 0.630000 1742.480000 1752.410000 ;
      RECT 1742.460000 0.000000 1742.480000 0.630000 ;
      RECT 1737.860000 0.000000 1742.040000 0.630000 ;
      RECT 1733.260000 0.000000 1737.440000 0.630000 ;
      RECT 1728.660000 0.000000 1732.840000 0.630000 ;
      RECT 1724.060000 0.000000 1728.240000 0.630000 ;
      RECT 1719.460000 0.000000 1723.640000 0.630000 ;
      RECT 1714.860000 0.000000 1719.040000 0.630000 ;
      RECT 1710.720000 0.000000 1714.440000 0.630000 ;
      RECT 1706.120000 0.000000 1710.300000 0.630000 ;
      RECT 1701.520000 0.000000 1705.700000 0.630000 ;
      RECT 1696.920000 0.000000 1701.100000 0.630000 ;
      RECT 1692.320000 0.000000 1696.500000 0.630000 ;
      RECT 1687.720000 0.000000 1691.900000 0.630000 ;
      RECT 1683.580000 0.000000 1687.300000 0.630000 ;
      RECT 1678.980000 0.000000 1683.160000 0.630000 ;
      RECT 1674.380000 0.000000 1678.560000 0.630000 ;
      RECT 1669.780000 0.000000 1673.960000 0.630000 ;
      RECT 1665.180000 0.000000 1669.360000 0.630000 ;
      RECT 1660.580000 0.000000 1664.760000 0.630000 ;
      RECT 1656.440000 0.000000 1660.160000 0.630000 ;
      RECT 1651.840000 0.000000 1656.020000 0.630000 ;
      RECT 1647.240000 0.000000 1651.420000 0.630000 ;
      RECT 1642.640000 0.000000 1646.820000 0.630000 ;
      RECT 1638.040000 0.000000 1642.220000 0.630000 ;
      RECT 1633.440000 0.000000 1637.620000 0.630000 ;
      RECT 1629.300000 0.000000 1633.020000 0.630000 ;
      RECT 1624.700000 0.000000 1628.880000 0.630000 ;
      RECT 1620.100000 0.000000 1624.280000 0.630000 ;
      RECT 1615.500000 0.000000 1619.680000 0.630000 ;
      RECT 1610.900000 0.000000 1615.080000 0.630000 ;
      RECT 1606.300000 0.000000 1610.480000 0.630000 ;
      RECT 1602.160000 0.000000 1605.880000 0.630000 ;
      RECT 1597.560000 0.000000 1601.740000 0.630000 ;
      RECT 1592.960000 0.000000 1597.140000 0.630000 ;
      RECT 1588.360000 0.000000 1592.540000 0.630000 ;
      RECT 1583.760000 0.000000 1587.940000 0.630000 ;
      RECT 1579.160000 0.000000 1583.340000 0.630000 ;
      RECT 1575.020000 0.000000 1578.740000 0.630000 ;
      RECT 1570.420000 0.000000 1574.600000 0.630000 ;
      RECT 1565.820000 0.000000 1570.000000 0.630000 ;
      RECT 1561.220000 0.000000 1565.400000 0.630000 ;
      RECT 1556.620000 0.000000 1560.800000 0.630000 ;
      RECT 1552.020000 0.000000 1556.200000 0.630000 ;
      RECT 1547.880000 0.000000 1551.600000 0.630000 ;
      RECT 1543.280000 0.000000 1547.460000 0.630000 ;
      RECT 1538.680000 0.000000 1542.860000 0.630000 ;
      RECT 1534.080000 0.000000 1538.260000 0.630000 ;
      RECT 1529.480000 0.000000 1533.660000 0.630000 ;
      RECT 1524.880000 0.000000 1529.060000 0.630000 ;
      RECT 1520.740000 0.000000 1524.460000 0.630000 ;
      RECT 1516.140000 0.000000 1520.320000 0.630000 ;
      RECT 1511.540000 0.000000 1515.720000 0.630000 ;
      RECT 1506.940000 0.000000 1511.120000 0.630000 ;
      RECT 1502.340000 0.000000 1506.520000 0.630000 ;
      RECT 1497.740000 0.000000 1501.920000 0.630000 ;
      RECT 1493.600000 0.000000 1497.320000 0.630000 ;
      RECT 1489.000000 0.000000 1493.180000 0.630000 ;
      RECT 1484.400000 0.000000 1488.580000 0.630000 ;
      RECT 1479.800000 0.000000 1483.980000 0.630000 ;
      RECT 1475.200000 0.000000 1479.380000 0.630000 ;
      RECT 1470.600000 0.000000 1474.780000 0.630000 ;
      RECT 1466.000000 0.000000 1470.180000 0.630000 ;
      RECT 1461.860000 0.000000 1465.580000 0.630000 ;
      RECT 1457.260000 0.000000 1461.440000 0.630000 ;
      RECT 1452.660000 0.000000 1456.840000 0.630000 ;
      RECT 1448.060000 0.000000 1452.240000 0.630000 ;
      RECT 1443.460000 0.000000 1447.640000 0.630000 ;
      RECT 1438.860000 0.000000 1443.040000 0.630000 ;
      RECT 1434.720000 0.000000 1438.440000 0.630000 ;
      RECT 1430.120000 0.000000 1434.300000 0.630000 ;
      RECT 1425.520000 0.000000 1429.700000 0.630000 ;
      RECT 1420.920000 0.000000 1425.100000 0.630000 ;
      RECT 1416.320000 0.000000 1420.500000 0.630000 ;
      RECT 1411.720000 0.000000 1415.900000 0.630000 ;
      RECT 1407.580000 0.000000 1411.300000 0.630000 ;
      RECT 1402.980000 0.000000 1407.160000 0.630000 ;
      RECT 1398.380000 0.000000 1402.560000 0.630000 ;
      RECT 1393.780000 0.000000 1397.960000 0.630000 ;
      RECT 1389.180000 0.000000 1393.360000 0.630000 ;
      RECT 1384.580000 0.000000 1388.760000 0.630000 ;
      RECT 1380.440000 0.000000 1384.160000 0.630000 ;
      RECT 1375.840000 0.000000 1380.020000 0.630000 ;
      RECT 1371.240000 0.000000 1375.420000 0.630000 ;
      RECT 1366.640000 0.000000 1370.820000 0.630000 ;
      RECT 1362.040000 0.000000 1366.220000 0.630000 ;
      RECT 1357.440000 0.000000 1361.620000 0.630000 ;
      RECT 1353.300000 0.000000 1357.020000 0.630000 ;
      RECT 1348.700000 0.000000 1352.880000 0.630000 ;
      RECT 1344.100000 0.000000 1348.280000 0.630000 ;
      RECT 1339.500000 0.000000 1343.680000 0.630000 ;
      RECT 1334.900000 0.000000 1339.080000 0.630000 ;
      RECT 1330.300000 0.000000 1334.480000 0.630000 ;
      RECT 1326.160000 0.000000 1329.880000 0.630000 ;
      RECT 1321.560000 0.000000 1325.740000 0.630000 ;
      RECT 1316.960000 0.000000 1321.140000 0.630000 ;
      RECT 1312.360000 0.000000 1316.540000 0.630000 ;
      RECT 1307.760000 0.000000 1311.940000 0.630000 ;
      RECT 1303.160000 0.000000 1307.340000 0.630000 ;
      RECT 1299.020000 0.000000 1302.740000 0.630000 ;
      RECT 1294.420000 0.000000 1298.600000 0.630000 ;
      RECT 1289.820000 0.000000 1294.000000 0.630000 ;
      RECT 1285.220000 0.000000 1289.400000 0.630000 ;
      RECT 1280.620000 0.000000 1284.800000 0.630000 ;
      RECT 1276.020000 0.000000 1280.200000 0.630000 ;
      RECT 1271.880000 0.000000 1275.600000 0.630000 ;
      RECT 1267.280000 0.000000 1271.460000 0.630000 ;
      RECT 1262.680000 0.000000 1266.860000 0.630000 ;
      RECT 1258.080000 0.000000 1262.260000 0.630000 ;
      RECT 1253.480000 0.000000 1257.660000 0.630000 ;
      RECT 1248.880000 0.000000 1253.060000 0.630000 ;
      RECT 1244.740000 0.000000 1248.460000 0.630000 ;
      RECT 1240.140000 0.000000 1244.320000 0.630000 ;
      RECT 1235.540000 0.000000 1239.720000 0.630000 ;
      RECT 1230.940000 0.000000 1235.120000 0.630000 ;
      RECT 1226.340000 0.000000 1230.520000 0.630000 ;
      RECT 1221.740000 0.000000 1225.920000 0.630000 ;
      RECT 1217.140000 0.000000 1221.320000 0.630000 ;
      RECT 1213.000000 0.000000 1216.720000 0.630000 ;
      RECT 1208.400000 0.000000 1212.580000 0.630000 ;
      RECT 1203.800000 0.000000 1207.980000 0.630000 ;
      RECT 1199.200000 0.000000 1203.380000 0.630000 ;
      RECT 1194.600000 0.000000 1198.780000 0.630000 ;
      RECT 1190.000000 0.000000 1194.180000 0.630000 ;
      RECT 1185.860000 0.000000 1189.580000 0.630000 ;
      RECT 1181.260000 0.000000 1185.440000 0.630000 ;
      RECT 1176.660000 0.000000 1180.840000 0.630000 ;
      RECT 1172.060000 0.000000 1176.240000 0.630000 ;
      RECT 1167.460000 0.000000 1171.640000 0.630000 ;
      RECT 1162.860000 0.000000 1167.040000 0.630000 ;
      RECT 1158.720000 0.000000 1162.440000 0.630000 ;
      RECT 1154.120000 0.000000 1158.300000 0.630000 ;
      RECT 1149.520000 0.000000 1153.700000 0.630000 ;
      RECT 1144.920000 0.000000 1149.100000 0.630000 ;
      RECT 1140.320000 0.000000 1144.500000 0.630000 ;
      RECT 1135.720000 0.000000 1139.900000 0.630000 ;
      RECT 1131.580000 0.000000 1135.300000 0.630000 ;
      RECT 1126.980000 0.000000 1131.160000 0.630000 ;
      RECT 1122.380000 0.000000 1126.560000 0.630000 ;
      RECT 1117.780000 0.000000 1121.960000 0.630000 ;
      RECT 1113.180000 0.000000 1117.360000 0.630000 ;
      RECT 1108.580000 0.000000 1112.760000 0.630000 ;
      RECT 1104.440000 0.000000 1108.160000 0.630000 ;
      RECT 1099.840000 0.000000 1104.020000 0.630000 ;
      RECT 1095.240000 0.000000 1099.420000 0.630000 ;
      RECT 1090.640000 0.000000 1094.820000 0.630000 ;
      RECT 1086.040000 0.000000 1090.220000 0.630000 ;
      RECT 1081.440000 0.000000 1085.620000 0.630000 ;
      RECT 1077.300000 0.000000 1081.020000 0.630000 ;
      RECT 1072.700000 0.000000 1076.880000 0.630000 ;
      RECT 1068.100000 0.000000 1072.280000 0.630000 ;
      RECT 1063.500000 0.000000 1067.680000 0.630000 ;
      RECT 1058.900000 0.000000 1063.080000 0.630000 ;
      RECT 1054.300000 0.000000 1058.480000 0.630000 ;
      RECT 1050.160000 0.000000 1053.880000 0.630000 ;
      RECT 1045.560000 0.000000 1049.740000 0.630000 ;
      RECT 1040.960000 0.000000 1045.140000 0.630000 ;
      RECT 1036.360000 0.000000 1040.540000 0.630000 ;
      RECT 1031.760000 0.000000 1035.940000 0.630000 ;
      RECT 1027.160000 0.000000 1031.340000 0.630000 ;
      RECT 1023.020000 0.000000 1026.740000 0.630000 ;
      RECT 1018.420000 0.000000 1022.600000 0.630000 ;
      RECT 1013.820000 0.000000 1018.000000 0.630000 ;
      RECT 1009.220000 0.000000 1013.400000 0.630000 ;
      RECT 1004.620000 0.000000 1008.800000 0.630000 ;
      RECT 1000.020000 0.000000 1004.200000 0.630000 ;
      RECT 995.420000 0.000000 999.600000 0.630000 ;
      RECT 991.280000 0.000000 995.000000 0.630000 ;
      RECT 986.680000 0.000000 990.860000 0.630000 ;
      RECT 982.080000 0.000000 986.260000 0.630000 ;
      RECT 977.480000 0.000000 981.660000 0.630000 ;
      RECT 972.880000 0.000000 977.060000 0.630000 ;
      RECT 968.280000 0.000000 972.460000 0.630000 ;
      RECT 964.140000 0.000000 967.860000 0.630000 ;
      RECT 959.540000 0.000000 963.720000 0.630000 ;
      RECT 954.940000 0.000000 959.120000 0.630000 ;
      RECT 950.340000 0.000000 954.520000 0.630000 ;
      RECT 945.740000 0.000000 949.920000 0.630000 ;
      RECT 941.140000 0.000000 945.320000 0.630000 ;
      RECT 937.000000 0.000000 940.720000 0.630000 ;
      RECT 932.400000 0.000000 936.580000 0.630000 ;
      RECT 927.800000 0.000000 931.980000 0.630000 ;
      RECT 923.200000 0.000000 927.380000 0.630000 ;
      RECT 918.600000 0.000000 922.780000 0.630000 ;
      RECT 914.000000 0.000000 918.180000 0.630000 ;
      RECT 909.860000 0.000000 913.580000 0.630000 ;
      RECT 905.260000 0.000000 909.440000 0.630000 ;
      RECT 900.660000 0.000000 904.840000 0.630000 ;
      RECT 896.060000 0.000000 900.240000 0.630000 ;
      RECT 891.460000 0.000000 895.640000 0.630000 ;
      RECT 886.860000 0.000000 891.040000 0.630000 ;
      RECT 882.720000 0.000000 886.440000 0.630000 ;
      RECT 878.120000 0.000000 882.300000 0.630000 ;
      RECT 873.520000 0.000000 877.700000 0.630000 ;
      RECT 868.920000 0.000000 873.100000 0.630000 ;
      RECT 864.320000 0.000000 868.500000 0.630000 ;
      RECT 859.720000 0.000000 863.900000 0.630000 ;
      RECT 855.580000 0.000000 859.300000 0.630000 ;
      RECT 850.980000 0.000000 855.160000 0.630000 ;
      RECT 846.380000 0.000000 850.560000 0.630000 ;
      RECT 841.780000 0.000000 845.960000 0.630000 ;
      RECT 837.180000 0.000000 841.360000 0.630000 ;
      RECT 832.580000 0.000000 836.760000 0.630000 ;
      RECT 828.440000 0.000000 832.160000 0.630000 ;
      RECT 823.840000 0.000000 828.020000 0.630000 ;
      RECT 819.240000 0.000000 823.420000 0.630000 ;
      RECT 814.640000 0.000000 818.820000 0.630000 ;
      RECT 810.040000 0.000000 814.220000 0.630000 ;
      RECT 805.440000 0.000000 809.620000 0.630000 ;
      RECT 801.300000 0.000000 805.020000 0.630000 ;
      RECT 796.700000 0.000000 800.880000 0.630000 ;
      RECT 792.100000 0.000000 796.280000 0.630000 ;
      RECT 787.500000 0.000000 791.680000 0.630000 ;
      RECT 782.900000 0.000000 787.080000 0.630000 ;
      RECT 778.300000 0.000000 782.480000 0.630000 ;
      RECT 774.160000 0.000000 777.880000 0.630000 ;
      RECT 769.560000 0.000000 773.740000 0.630000 ;
      RECT 764.960000 0.000000 769.140000 0.630000 ;
      RECT 760.360000 0.000000 764.540000 0.630000 ;
      RECT 755.760000 0.000000 759.940000 0.630000 ;
      RECT 751.160000 0.000000 755.340000 0.630000 ;
      RECT 746.560000 0.000000 750.740000 0.630000 ;
      RECT 742.420000 0.000000 746.140000 0.630000 ;
      RECT 737.820000 0.000000 742.000000 0.630000 ;
      RECT 733.220000 0.000000 737.400000 0.630000 ;
      RECT 728.620000 0.000000 732.800000 0.630000 ;
      RECT 724.020000 0.000000 728.200000 0.630000 ;
      RECT 719.420000 0.000000 723.600000 0.630000 ;
      RECT 715.280000 0.000000 719.000000 0.630000 ;
      RECT 710.680000 0.000000 714.860000 0.630000 ;
      RECT 706.080000 0.000000 710.260000 0.630000 ;
      RECT 701.480000 0.000000 705.660000 0.630000 ;
      RECT 696.880000 0.000000 701.060000 0.630000 ;
      RECT 692.280000 0.000000 696.460000 0.630000 ;
      RECT 688.140000 0.000000 691.860000 0.630000 ;
      RECT 683.540000 0.000000 687.720000 0.630000 ;
      RECT 678.940000 0.000000 683.120000 0.630000 ;
      RECT 674.340000 0.000000 678.520000 0.630000 ;
      RECT 669.740000 0.000000 673.920000 0.630000 ;
      RECT 665.140000 0.000000 669.320000 0.630000 ;
      RECT 661.000000 0.000000 664.720000 0.630000 ;
      RECT 656.400000 0.000000 660.580000 0.630000 ;
      RECT 651.800000 0.000000 655.980000 0.630000 ;
      RECT 647.200000 0.000000 651.380000 0.630000 ;
      RECT 642.600000 0.000000 646.780000 0.630000 ;
      RECT 638.000000 0.000000 642.180000 0.630000 ;
      RECT 633.860000 0.000000 637.580000 0.630000 ;
      RECT 629.260000 0.000000 633.440000 0.630000 ;
      RECT 624.660000 0.000000 628.840000 0.630000 ;
      RECT 620.060000 0.000000 624.240000 0.630000 ;
      RECT 615.460000 0.000000 619.640000 0.630000 ;
      RECT 610.860000 0.000000 615.040000 0.630000 ;
      RECT 606.720000 0.000000 610.440000 0.630000 ;
      RECT 602.120000 0.000000 606.300000 0.630000 ;
      RECT 597.520000 0.000000 601.700000 0.630000 ;
      RECT 592.920000 0.000000 597.100000 0.630000 ;
      RECT 588.320000 0.000000 592.500000 0.630000 ;
      RECT 583.720000 0.000000 587.900000 0.630000 ;
      RECT 579.580000 0.000000 583.300000 0.630000 ;
      RECT 574.980000 0.000000 579.160000 0.630000 ;
      RECT 570.380000 0.000000 574.560000 0.630000 ;
      RECT 565.780000 0.000000 569.960000 0.630000 ;
      RECT 561.180000 0.000000 565.360000 0.630000 ;
      RECT 556.580000 0.000000 560.760000 0.630000 ;
      RECT 552.440000 0.000000 556.160000 0.630000 ;
      RECT 547.840000 0.000000 552.020000 0.630000 ;
      RECT 543.240000 0.000000 547.420000 0.630000 ;
      RECT 538.640000 0.000000 542.820000 0.630000 ;
      RECT 534.040000 0.000000 538.220000 0.630000 ;
      RECT 529.440000 0.000000 533.620000 0.630000 ;
      RECT 525.300000 0.000000 529.020000 0.630000 ;
      RECT 520.700000 0.000000 524.880000 0.630000 ;
      RECT 516.100000 0.000000 520.280000 0.630000 ;
      RECT 511.500000 0.000000 515.680000 0.630000 ;
      RECT 506.900000 0.000000 511.080000 0.630000 ;
      RECT 502.300000 0.000000 506.480000 0.630000 ;
      RECT 498.160000 0.000000 501.880000 0.630000 ;
      RECT 493.560000 0.000000 497.740000 0.630000 ;
      RECT 488.960000 0.000000 493.140000 0.630000 ;
      RECT 484.360000 0.000000 488.540000 0.630000 ;
      RECT 479.760000 0.000000 483.940000 0.630000 ;
      RECT 475.160000 0.000000 479.340000 0.630000 ;
      RECT 470.560000 0.000000 474.740000 0.630000 ;
      RECT 466.420000 0.000000 470.140000 0.630000 ;
      RECT 461.820000 0.000000 466.000000 0.630000 ;
      RECT 457.220000 0.000000 461.400000 0.630000 ;
      RECT 452.620000 0.000000 456.800000 0.630000 ;
      RECT 448.020000 0.000000 452.200000 0.630000 ;
      RECT 443.420000 0.000000 447.600000 0.630000 ;
      RECT 439.280000 0.000000 443.000000 0.630000 ;
      RECT 434.680000 0.000000 438.860000 0.630000 ;
      RECT 430.080000 0.000000 434.260000 0.630000 ;
      RECT 425.480000 0.000000 429.660000 0.630000 ;
      RECT 420.880000 0.000000 425.060000 0.630000 ;
      RECT 416.280000 0.000000 420.460000 0.630000 ;
      RECT 412.140000 0.000000 415.860000 0.630000 ;
      RECT 407.540000 0.000000 411.720000 0.630000 ;
      RECT 402.940000 0.000000 407.120000 0.630000 ;
      RECT 398.340000 0.000000 402.520000 0.630000 ;
      RECT 393.740000 0.000000 397.920000 0.630000 ;
      RECT 389.140000 0.000000 393.320000 0.630000 ;
      RECT 385.000000 0.000000 388.720000 0.630000 ;
      RECT 380.400000 0.000000 384.580000 0.630000 ;
      RECT 375.800000 0.000000 379.980000 0.630000 ;
      RECT 371.200000 0.000000 375.380000 0.630000 ;
      RECT 366.600000 0.000000 370.780000 0.630000 ;
      RECT 362.000000 0.000000 366.180000 0.630000 ;
      RECT 357.860000 0.000000 361.580000 0.630000 ;
      RECT 353.260000 0.000000 357.440000 0.630000 ;
      RECT 348.660000 0.000000 352.840000 0.630000 ;
      RECT 344.060000 0.000000 348.240000 0.630000 ;
      RECT 339.460000 0.000000 343.640000 0.630000 ;
      RECT 334.860000 0.000000 339.040000 0.630000 ;
      RECT 330.720000 0.000000 334.440000 0.630000 ;
      RECT 326.120000 0.000000 330.300000 0.630000 ;
      RECT 321.520000 0.000000 325.700000 0.630000 ;
      RECT 316.920000 0.000000 321.100000 0.630000 ;
      RECT 312.320000 0.000000 316.500000 0.630000 ;
      RECT 307.720000 0.000000 311.900000 0.630000 ;
      RECT 303.580000 0.000000 307.300000 0.630000 ;
      RECT 298.980000 0.000000 303.160000 0.630000 ;
      RECT 294.380000 0.000000 298.560000 0.630000 ;
      RECT 289.780000 0.000000 293.960000 0.630000 ;
      RECT 285.180000 0.000000 289.360000 0.630000 ;
      RECT 280.580000 0.000000 284.760000 0.630000 ;
      RECT 276.440000 0.000000 280.160000 0.630000 ;
      RECT 271.840000 0.000000 276.020000 0.630000 ;
      RECT 267.240000 0.000000 271.420000 0.630000 ;
      RECT 262.640000 0.000000 266.820000 0.630000 ;
      RECT 258.040000 0.000000 262.220000 0.630000 ;
      RECT 253.440000 0.000000 257.620000 0.630000 ;
      RECT 248.840000 0.000000 253.020000 0.630000 ;
      RECT 244.700000 0.000000 248.420000 0.630000 ;
      RECT 240.100000 0.000000 244.280000 0.630000 ;
      RECT 235.500000 0.000000 239.680000 0.630000 ;
      RECT 230.900000 0.000000 235.080000 0.630000 ;
      RECT 226.300000 0.000000 230.480000 0.630000 ;
      RECT 221.700000 0.000000 225.880000 0.630000 ;
      RECT 217.560000 0.000000 221.280000 0.630000 ;
      RECT 212.960000 0.000000 217.140000 0.630000 ;
      RECT 208.360000 0.000000 212.540000 0.630000 ;
      RECT 203.760000 0.000000 207.940000 0.630000 ;
      RECT 199.160000 0.000000 203.340000 0.630000 ;
      RECT 194.560000 0.000000 198.740000 0.630000 ;
      RECT 190.420000 0.000000 194.140000 0.630000 ;
      RECT 185.820000 0.000000 190.000000 0.630000 ;
      RECT 181.220000 0.000000 185.400000 0.630000 ;
      RECT 176.620000 0.000000 180.800000 0.630000 ;
      RECT 172.020000 0.000000 176.200000 0.630000 ;
      RECT 167.420000 0.000000 171.600000 0.630000 ;
      RECT 163.280000 0.000000 167.000000 0.630000 ;
      RECT 158.680000 0.000000 162.860000 0.630000 ;
      RECT 154.080000 0.000000 158.260000 0.630000 ;
      RECT 149.480000 0.000000 153.660000 0.630000 ;
      RECT 144.880000 0.000000 149.060000 0.630000 ;
      RECT 140.280000 0.000000 144.460000 0.630000 ;
      RECT 136.140000 0.000000 139.860000 0.630000 ;
      RECT 131.540000 0.000000 135.720000 0.630000 ;
      RECT 126.940000 0.000000 131.120000 0.630000 ;
      RECT 122.340000 0.000000 126.520000 0.630000 ;
      RECT 117.740000 0.000000 121.920000 0.630000 ;
      RECT 113.140000 0.000000 117.320000 0.630000 ;
      RECT 109.000000 0.000000 112.720000 0.630000 ;
      RECT 104.400000 0.000000 108.580000 0.630000 ;
      RECT 99.800000 0.000000 103.980000 0.630000 ;
      RECT 95.200000 0.000000 99.380000 0.630000 ;
      RECT 90.600000 0.000000 94.780000 0.630000 ;
      RECT 86.000000 0.000000 90.180000 0.630000 ;
      RECT 81.860000 0.000000 85.580000 0.630000 ;
      RECT 77.260000 0.000000 81.440000 0.630000 ;
      RECT 72.660000 0.000000 76.840000 0.630000 ;
      RECT 68.060000 0.000000 72.240000 0.630000 ;
      RECT 63.460000 0.000000 67.640000 0.630000 ;
      RECT 58.860000 0.000000 63.040000 0.630000 ;
      RECT 54.720000 0.000000 58.440000 0.630000 ;
      RECT 50.120000 0.000000 54.300000 0.630000 ;
      RECT 45.520000 0.000000 49.700000 0.630000 ;
      RECT 40.920000 0.000000 45.100000 0.630000 ;
      RECT 36.320000 0.000000 40.500000 0.630000 ;
      RECT 31.720000 0.000000 35.900000 0.630000 ;
      RECT 27.580000 0.000000 31.300000 0.630000 ;
      RECT 22.980000 0.000000 27.160000 0.630000 ;
      RECT 18.380000 0.000000 22.560000 0.630000 ;
      RECT 13.780000 0.000000 17.960000 0.630000 ;
      RECT 9.180000 0.000000 13.360000 0.630000 ;
      RECT 4.580000 0.000000 8.760000 0.630000 ;
      RECT 0.440000 0.000000 4.160000 0.630000 ;
      RECT 0.000000 0.000000 0.020000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 1752.470000 1741.380000 1753.040000 ;
      RECT 1.100000 1752.180000 1741.380000 1752.470000 ;
      RECT 1.100000 1751.570000 1742.480000 1752.180000 ;
      RECT 0.000000 1712.820000 1742.480000 1751.570000 ;
      RECT 0.000000 1711.920000 1741.380000 1712.820000 ;
      RECT 0.000000 1709.770000 1742.480000 1711.920000 ;
      RECT 1.100000 1708.870000 1742.480000 1709.770000 ;
      RECT 0.000000 1673.170000 1742.480000 1708.870000 ;
      RECT 0.000000 1672.270000 1741.380000 1673.170000 ;
      RECT 0.000000 1667.070000 1742.480000 1672.270000 ;
      RECT 1.100000 1666.170000 1742.480000 1667.070000 ;
      RECT 0.000000 1633.520000 1742.480000 1666.170000 ;
      RECT 0.000000 1632.620000 1741.380000 1633.520000 ;
      RECT 0.000000 1624.370000 1742.480000 1632.620000 ;
      RECT 1.100000 1623.470000 1742.480000 1624.370000 ;
      RECT 0.000000 1593.260000 1742.480000 1623.470000 ;
      RECT 0.000000 1592.360000 1741.380000 1593.260000 ;
      RECT 0.000000 1581.670000 1742.480000 1592.360000 ;
      RECT 1.100000 1580.770000 1742.480000 1581.670000 ;
      RECT 0.000000 1553.610000 1742.480000 1580.770000 ;
      RECT 0.000000 1552.710000 1741.380000 1553.610000 ;
      RECT 0.000000 1538.970000 1742.480000 1552.710000 ;
      RECT 1.100000 1538.070000 1742.480000 1538.970000 ;
      RECT 0.000000 1513.960000 1742.480000 1538.070000 ;
      RECT 0.000000 1513.060000 1741.380000 1513.960000 ;
      RECT 0.000000 1496.270000 1742.480000 1513.060000 ;
      RECT 1.100000 1495.370000 1742.480000 1496.270000 ;
      RECT 0.000000 1474.310000 1742.480000 1495.370000 ;
      RECT 0.000000 1473.410000 1741.380000 1474.310000 ;
      RECT 0.000000 1453.570000 1742.480000 1473.410000 ;
      RECT 1.100000 1452.670000 1742.480000 1453.570000 ;
      RECT 0.000000 1434.050000 1742.480000 1452.670000 ;
      RECT 0.000000 1433.150000 1741.380000 1434.050000 ;
      RECT 0.000000 1410.870000 1742.480000 1433.150000 ;
      RECT 1.100000 1409.970000 1742.480000 1410.870000 ;
      RECT 0.000000 1394.400000 1742.480000 1409.970000 ;
      RECT 0.000000 1393.500000 1741.380000 1394.400000 ;
      RECT 0.000000 1368.170000 1742.480000 1393.500000 ;
      RECT 1.100000 1367.270000 1742.480000 1368.170000 ;
      RECT 0.000000 1354.750000 1742.480000 1367.270000 ;
      RECT 0.000000 1353.850000 1741.380000 1354.750000 ;
      RECT 0.000000 1325.470000 1742.480000 1353.850000 ;
      RECT 1.100000 1324.570000 1742.480000 1325.470000 ;
      RECT 0.000000 1315.100000 1742.480000 1324.570000 ;
      RECT 0.000000 1314.200000 1741.380000 1315.100000 ;
      RECT 0.000000 1282.770000 1742.480000 1314.200000 ;
      RECT 1.100000 1281.870000 1742.480000 1282.770000 ;
      RECT 0.000000 1274.840000 1742.480000 1281.870000 ;
      RECT 0.000000 1273.940000 1741.380000 1274.840000 ;
      RECT 0.000000 1240.070000 1742.480000 1273.940000 ;
      RECT 1.100000 1239.170000 1742.480000 1240.070000 ;
      RECT 0.000000 1235.190000 1742.480000 1239.170000 ;
      RECT 0.000000 1234.290000 1741.380000 1235.190000 ;
      RECT 0.000000 1197.370000 1742.480000 1234.290000 ;
      RECT 1.100000 1196.470000 1742.480000 1197.370000 ;
      RECT 0.000000 1195.540000 1742.480000 1196.470000 ;
      RECT 0.000000 1194.640000 1741.380000 1195.540000 ;
      RECT 0.000000 1155.280000 1742.480000 1194.640000 ;
      RECT 0.000000 1154.670000 1741.380000 1155.280000 ;
      RECT 1.100000 1154.380000 1741.380000 1154.670000 ;
      RECT 1.100000 1153.770000 1742.480000 1154.380000 ;
      RECT 0.000000 1115.630000 1742.480000 1153.770000 ;
      RECT 0.000000 1114.730000 1741.380000 1115.630000 ;
      RECT 0.000000 1111.970000 1742.480000 1114.730000 ;
      RECT 1.100000 1111.070000 1742.480000 1111.970000 ;
      RECT 0.000000 1075.980000 1742.480000 1111.070000 ;
      RECT 0.000000 1075.080000 1741.380000 1075.980000 ;
      RECT 0.000000 1069.270000 1742.480000 1075.080000 ;
      RECT 1.100000 1068.370000 1742.480000 1069.270000 ;
      RECT 0.000000 1036.330000 1742.480000 1068.370000 ;
      RECT 0.000000 1035.430000 1741.380000 1036.330000 ;
      RECT 0.000000 1026.570000 1742.480000 1035.430000 ;
      RECT 1.100000 1025.670000 1742.480000 1026.570000 ;
      RECT 0.000000 996.070000 1742.480000 1025.670000 ;
      RECT 0.000000 995.170000 1741.380000 996.070000 ;
      RECT 0.000000 983.870000 1742.480000 995.170000 ;
      RECT 1.100000 982.970000 1742.480000 983.870000 ;
      RECT 0.000000 956.420000 1742.480000 982.970000 ;
      RECT 0.000000 955.520000 1741.380000 956.420000 ;
      RECT 0.000000 941.170000 1742.480000 955.520000 ;
      RECT 1.100000 940.270000 1742.480000 941.170000 ;
      RECT 0.000000 916.770000 1742.480000 940.270000 ;
      RECT 0.000000 915.870000 1741.380000 916.770000 ;
      RECT 0.000000 898.470000 1742.480000 915.870000 ;
      RECT 1.100000 897.570000 1742.480000 898.470000 ;
      RECT 0.000000 876.510000 1742.480000 897.570000 ;
      RECT 0.000000 875.610000 1741.380000 876.510000 ;
      RECT 0.000000 855.160000 1742.480000 875.610000 ;
      RECT 1.100000 854.260000 1742.480000 855.160000 ;
      RECT 0.000000 836.860000 1742.480000 854.260000 ;
      RECT 0.000000 835.960000 1741.380000 836.860000 ;
      RECT 0.000000 812.460000 1742.480000 835.960000 ;
      RECT 1.100000 811.560000 1742.480000 812.460000 ;
      RECT 0.000000 797.210000 1742.480000 811.560000 ;
      RECT 0.000000 796.310000 1741.380000 797.210000 ;
      RECT 0.000000 769.760000 1742.480000 796.310000 ;
      RECT 1.100000 768.860000 1742.480000 769.760000 ;
      RECT 0.000000 757.560000 1742.480000 768.860000 ;
      RECT 0.000000 756.660000 1741.380000 757.560000 ;
      RECT 0.000000 727.060000 1742.480000 756.660000 ;
      RECT 1.100000 726.160000 1742.480000 727.060000 ;
      RECT 0.000000 717.300000 1742.480000 726.160000 ;
      RECT 0.000000 716.400000 1741.380000 717.300000 ;
      RECT 0.000000 684.360000 1742.480000 716.400000 ;
      RECT 1.100000 683.460000 1742.480000 684.360000 ;
      RECT 0.000000 677.650000 1742.480000 683.460000 ;
      RECT 0.000000 676.750000 1741.380000 677.650000 ;
      RECT 0.000000 641.660000 1742.480000 676.750000 ;
      RECT 1.100000 640.760000 1742.480000 641.660000 ;
      RECT 0.000000 638.000000 1742.480000 640.760000 ;
      RECT 0.000000 637.100000 1741.380000 638.000000 ;
      RECT 0.000000 598.960000 1742.480000 637.100000 ;
      RECT 1.100000 598.350000 1742.480000 598.960000 ;
      RECT 1.100000 598.060000 1741.380000 598.350000 ;
      RECT 0.000000 597.450000 1741.380000 598.060000 ;
      RECT 0.000000 558.090000 1742.480000 597.450000 ;
      RECT 0.000000 557.190000 1741.380000 558.090000 ;
      RECT 0.000000 556.260000 1742.480000 557.190000 ;
      RECT 1.100000 555.360000 1742.480000 556.260000 ;
      RECT 0.000000 518.440000 1742.480000 555.360000 ;
      RECT 0.000000 517.540000 1741.380000 518.440000 ;
      RECT 0.000000 513.560000 1742.480000 517.540000 ;
      RECT 1.100000 512.660000 1742.480000 513.560000 ;
      RECT 0.000000 478.790000 1742.480000 512.660000 ;
      RECT 0.000000 477.890000 1741.380000 478.790000 ;
      RECT 0.000000 470.860000 1742.480000 477.890000 ;
      RECT 1.100000 469.960000 1742.480000 470.860000 ;
      RECT 0.000000 438.530000 1742.480000 469.960000 ;
      RECT 0.000000 437.630000 1741.380000 438.530000 ;
      RECT 0.000000 428.160000 1742.480000 437.630000 ;
      RECT 1.100000 427.260000 1742.480000 428.160000 ;
      RECT 0.000000 398.880000 1742.480000 427.260000 ;
      RECT 0.000000 397.980000 1741.380000 398.880000 ;
      RECT 0.000000 385.460000 1742.480000 397.980000 ;
      RECT 1.100000 384.560000 1742.480000 385.460000 ;
      RECT 0.000000 359.230000 1742.480000 384.560000 ;
      RECT 0.000000 358.330000 1741.380000 359.230000 ;
      RECT 0.000000 342.760000 1742.480000 358.330000 ;
      RECT 1.100000 341.860000 1742.480000 342.760000 ;
      RECT 0.000000 319.580000 1742.480000 341.860000 ;
      RECT 0.000000 318.680000 1741.380000 319.580000 ;
      RECT 0.000000 300.060000 1742.480000 318.680000 ;
      RECT 1.100000 299.160000 1742.480000 300.060000 ;
      RECT 0.000000 279.320000 1742.480000 299.160000 ;
      RECT 0.000000 278.420000 1741.380000 279.320000 ;
      RECT 0.000000 257.360000 1742.480000 278.420000 ;
      RECT 1.100000 256.460000 1742.480000 257.360000 ;
      RECT 0.000000 239.670000 1742.480000 256.460000 ;
      RECT 0.000000 238.770000 1741.380000 239.670000 ;
      RECT 0.000000 214.660000 1742.480000 238.770000 ;
      RECT 1.100000 213.760000 1742.480000 214.660000 ;
      RECT 0.000000 200.020000 1742.480000 213.760000 ;
      RECT 0.000000 199.120000 1741.380000 200.020000 ;
      RECT 0.000000 171.960000 1742.480000 199.120000 ;
      RECT 1.100000 171.060000 1742.480000 171.960000 ;
      RECT 0.000000 160.370000 1742.480000 171.060000 ;
      RECT 0.000000 159.470000 1741.380000 160.370000 ;
      RECT 0.000000 129.260000 1742.480000 159.470000 ;
      RECT 1.100000 128.360000 1742.480000 129.260000 ;
      RECT 0.000000 120.110000 1742.480000 128.360000 ;
      RECT 0.000000 119.210000 1741.380000 120.110000 ;
      RECT 0.000000 86.560000 1742.480000 119.210000 ;
      RECT 1.100000 85.660000 1742.480000 86.560000 ;
      RECT 0.000000 80.460000 1742.480000 85.660000 ;
      RECT 0.000000 79.560000 1741.380000 80.460000 ;
      RECT 0.000000 43.860000 1742.480000 79.560000 ;
      RECT 1.100000 42.960000 1742.480000 43.860000 ;
      RECT 0.000000 40.810000 1742.480000 42.960000 ;
      RECT 0.000000 39.910000 1741.380000 40.810000 ;
      RECT 0.000000 1.160000 1742.480000 39.910000 ;
      RECT 1.100000 0.260000 1741.380000 1.160000 ;
      RECT 0.000000 0.000000 1742.480000 0.260000 ;
    LAYER met4 ;
      RECT 0.000000 1748.290000 1742.480000 1753.040000 ;
      RECT 9.390000 1741.490000 1733.090000 1748.290000 ;
      RECT 1732.090000 10.530000 1733.090000 1741.490000 ;
      RECT 16.190000 10.530000 1726.290000 1741.490000 ;
      RECT 9.390000 10.530000 10.390000 1741.490000 ;
      RECT 1738.890000 3.730000 1742.480000 1748.290000 ;
      RECT 9.390000 3.730000 1733.090000 10.530000 ;
      RECT 0.000000 3.730000 3.590000 1748.290000 ;
      RECT 0.000000 0.000000 1742.480000 3.730000 ;
  END
END Ibtida_top_dffram_cv

END LIBRARY
